module inv(in, out);
input in;
output out;
assign out = ~in;
endmodule

module nand2(a, b, out);
input a, b;
output out;
assign out = ~(a & b);
endmodule

module nand3(a, b, c, out);
input a, b, c;
output out;
assign out = ~(a & b & c);
endmodule

module nand4(a, b, c, d, out);
input a, b, c, d;
output out;
assign out = ~(a & b & c & d);
endmodule

module nor2(a, b, out);
input a, b;
output out;
assign out = ~(a | b);
endmodule

module nor3(a, b, c, out);
input a, b, c;
output out;
assign out = ~(a | b | c);
endmodule

module xor2(a, b, out);
input a, b;
output out;
assign out = (a ^ b);
endmodule

module aoi12(a, b, c, out);
input a, b, c;
output out;
assign out = ~(a | (b & c));
endmodule

module aoi22(a, b, c, d, out);
input a, b, c, d;
output out;
assign out = ~((a & b) | (c & d));
endmodule

module oai12(a, b, c, out);
input a, b, c;
output out;
assign out = ~(a & (b | c));
endmodule

module oai22(a, b, c, d, out);
input a, b, c, d;
output out;
assign out = ~((a | b) & (c | d));
endmodule

module dff( d, gclk, rnot, q);
input d, gclk, rnot;
output q;
reg q;
always @(posedge gclk or negedge rnot)
  if (rnot == 1'b0)
    q = 1'b0;
  else
    q = d;
endmodule


/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : O-2018.06-SP1
// Date      : Sat Oct 28 11:55:25 2023
/////////////////////////////////////////////////////////////


module matrix_alu_mapped ( clk, resetn, A, B, op, C );
  input [31:0] A;
  input [31:0] B;
  input [1:0] op;
  output [127:0] C;
  input clk, resetn;
  wire   N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33,
         N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47,
         N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61,
         N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75,
         N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89,
         N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102,
         N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113,
         N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124,
         N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135,
         N136, N137, N139, N140, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[0] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[3] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[5] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[7] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[0] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[7] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[0] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[3] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[5] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[7] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[0] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[7] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[0] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[3] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[5] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[7] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[0] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[7] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[0] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[3] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[5] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[7] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[0] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ,
         \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[7] ,
         \mat_kron/mult_40/FS_1/P[0][0][1] ,
         \mat_kron/mult_40/FS_1/P[0][0][2] ,
         \mat_kron/mult_40/FS_1/P[0][0][3] ,
         \mat_kron/mult_40/FS_1/P[0][1][1] ,
         \mat_kron/mult_40/FS_1/TEMP_P[0][0][0] ,
         \mat_kron/mult_40/FS_1/TEMP_P[0][1][0] , \mat_kron/mult_40/A1[0] ,
         \mat_kron/mult_40/A1[1] , \mat_kron/mult_40/A1[2] ,
         \mat_kron/mult_40/A1[3] , \mat_kron/mult_40/A1[4] ,
         \mat_kron/mult_40/A1[5] , \mat_kron/mult_40/A_notx[0] ,
         \mat_kron/mult_40/B_notx[0] , \mat_kron/mult_40/ab[0][1] ,
         \mat_kron/mult_40/ab[0][2] , \mat_kron/mult_40/ab[0][3] ,
         \mat_kron/mult_40/ab[0][4] , \mat_kron/mult_40/ab[0][5] ,
         \mat_kron/mult_40/ab[0][6] , \mat_kron/mult_40/ab[0][7] ,
         \mat_kron/mult_40/ab[1][0] , \mat_kron/mult_40/ab[1][1] ,
         \mat_kron/mult_40/ab[1][2] , \mat_kron/mult_40/ab[1][3] ,
         \mat_kron/mult_40/ab[1][4] , \mat_kron/mult_40/ab[1][5] ,
         \mat_kron/mult_40/ab[1][6] , \mat_kron/mult_40/ab[2][0] ,
         \mat_kron/mult_40/ab[2][1] , \mat_kron/mult_40/ab[2][2] ,
         \mat_kron/mult_40/ab[2][3] , \mat_kron/mult_40/ab[2][4] ,
         \mat_kron/mult_40/ab[2][5] , \mat_kron/mult_40/ab[3][0] ,
         \mat_kron/mult_40/ab[3][1] , \mat_kron/mult_40/ab[3][2] ,
         \mat_kron/mult_40/ab[3][3] , \mat_kron/mult_40/ab[3][4] ,
         \mat_kron/mult_40/ab[4][0] , \mat_kron/mult_40/ab[4][1] ,
         \mat_kron/mult_40/ab[4][2] , \mat_kron/mult_40/ab[4][3] ,
         \mat_kron/mult_40/ab[5][0] , \mat_kron/mult_40/ab[5][1] ,
         \mat_kron/mult_40/ab[5][2] , \mat_kron/mult_40/ab[6][0] ,
         \mat_kron/mult_40/ab[6][1] , \mat_kron/mult_40/ab[7][0] ,
         \mat_kron/mult_40_G2_G1_G1_G1/FS_1/P[0][0][1] ,
         \mat_kron/mult_40_G2_G1_G1_G1/FS_1/P[0][0][2] ,
         \mat_kron/mult_40_G2_G1_G1_G1/FS_1/P[0][0][3] ,
         \mat_kron/mult_40_G2_G1_G1_G1/FS_1/P[0][1][1] ,
         \mat_kron/mult_40_G2_G1_G1_G1/FS_1/TEMP_P[0][0][0] ,
         \mat_kron/mult_40_G2_G1_G1_G1/FS_1/TEMP_P[0][1][0] ,
         \mat_kron/mult_40_G2_G1_G1_G1/A1[0] ,
         \mat_kron/mult_40_G2_G1_G1_G1/A1[1] ,
         \mat_kron/mult_40_G2_G1_G1_G1/A1[2] ,
         \mat_kron/mult_40_G2_G1_G1_G1/A1[3] ,
         \mat_kron/mult_40_G2_G1_G1_G1/A1[4] ,
         \mat_kron/mult_40_G2_G1_G1_G1/A1[5] ,
         \mat_kron/mult_40_G2_G1_G1_G1/A_notx[0] ,
         \mat_kron/mult_40_G2_G1_G1_G1/B_notx[0] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[0][1] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[0][2] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[0][3] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[0][4] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[0][5] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[0][6] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[0][7] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[1][0] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[1][1] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[1][2] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[1][3] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[1][4] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[1][5] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[1][6] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[2][0] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[2][1] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[2][2] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[2][3] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[2][4] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[2][5] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[3][0] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[3][1] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[3][2] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[3][3] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[3][4] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[4][0] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[4][1] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[4][2] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[4][3] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[5][0] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[5][1] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[5][2] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[6][0] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[6][1] ,
         \mat_kron/mult_40_G2_G1_G1_G1/ab[7][0] ,
         \mat_kron/mult_40_G2_G1_G1/FS_1/P[0][0][1] ,
         \mat_kron/mult_40_G2_G1_G1/FS_1/P[0][0][2] ,
         \mat_kron/mult_40_G2_G1_G1/FS_1/P[0][0][3] ,
         \mat_kron/mult_40_G2_G1_G1/FS_1/P[0][1][1] ,
         \mat_kron/mult_40_G2_G1_G1/FS_1/TEMP_P[0][0][0] ,
         \mat_kron/mult_40_G2_G1_G1/FS_1/TEMP_P[0][1][0] ,
         \mat_kron/mult_40_G2_G1_G1/A1[0] , \mat_kron/mult_40_G2_G1_G1/A1[1] ,
         \mat_kron/mult_40_G2_G1_G1/A1[2] , \mat_kron/mult_40_G2_G1_G1/A1[3] ,
         \mat_kron/mult_40_G2_G1_G1/A1[4] , \mat_kron/mult_40_G2_G1_G1/A1[5] ,
         \mat_kron/mult_40_G2_G1_G1/A_notx[0] ,
         \mat_kron/mult_40_G2_G1_G1/B_notx[0] ,
         \mat_kron/mult_40_G2_G1_G1/ab[0][1] ,
         \mat_kron/mult_40_G2_G1_G1/ab[0][2] ,
         \mat_kron/mult_40_G2_G1_G1/ab[0][3] ,
         \mat_kron/mult_40_G2_G1_G1/ab[0][4] ,
         \mat_kron/mult_40_G2_G1_G1/ab[0][5] ,
         \mat_kron/mult_40_G2_G1_G1/ab[0][6] ,
         \mat_kron/mult_40_G2_G1_G1/ab[0][7] ,
         \mat_kron/mult_40_G2_G1_G1/ab[1][0] ,
         \mat_kron/mult_40_G2_G1_G1/ab[1][1] ,
         \mat_kron/mult_40_G2_G1_G1/ab[1][2] ,
         \mat_kron/mult_40_G2_G1_G1/ab[1][3] ,
         \mat_kron/mult_40_G2_G1_G1/ab[1][4] ,
         \mat_kron/mult_40_G2_G1_G1/ab[1][5] ,
         \mat_kron/mult_40_G2_G1_G1/ab[1][6] ,
         \mat_kron/mult_40_G2_G1_G1/ab[2][0] ,
         \mat_kron/mult_40_G2_G1_G1/ab[2][1] ,
         \mat_kron/mult_40_G2_G1_G1/ab[2][2] ,
         \mat_kron/mult_40_G2_G1_G1/ab[2][3] ,
         \mat_kron/mult_40_G2_G1_G1/ab[2][4] ,
         \mat_kron/mult_40_G2_G1_G1/ab[2][5] ,
         \mat_kron/mult_40_G2_G1_G1/ab[3][0] ,
         \mat_kron/mult_40_G2_G1_G1/ab[3][1] ,
         \mat_kron/mult_40_G2_G1_G1/ab[3][2] ,
         \mat_kron/mult_40_G2_G1_G1/ab[3][3] ,
         \mat_kron/mult_40_G2_G1_G1/ab[3][4] ,
         \mat_kron/mult_40_G2_G1_G1/ab[4][0] ,
         \mat_kron/mult_40_G2_G1_G1/ab[4][1] ,
         \mat_kron/mult_40_G2_G1_G1/ab[4][2] ,
         \mat_kron/mult_40_G2_G1_G1/ab[4][3] ,
         \mat_kron/mult_40_G2_G1_G1/ab[5][0] ,
         \mat_kron/mult_40_G2_G1_G1/ab[5][1] ,
         \mat_kron/mult_40_G2_G1_G1/ab[5][2] ,
         \mat_kron/mult_40_G2_G1_G1/ab[6][0] ,
         \mat_kron/mult_40_G2_G1_G1/ab[6][1] ,
         \mat_kron/mult_40_G2_G1_G1/ab[7][0] ,
         \mat_kron/mult_40_G2_G2_G1_G1/FS_1/P[0][0][1] ,
         \mat_kron/mult_40_G2_G2_G1_G1/FS_1/P[0][0][2] ,
         \mat_kron/mult_40_G2_G2_G1_G1/FS_1/P[0][0][3] ,
         \mat_kron/mult_40_G2_G2_G1_G1/FS_1/P[0][1][1] ,
         \mat_kron/mult_40_G2_G2_G1_G1/FS_1/TEMP_P[0][0][0] ,
         \mat_kron/mult_40_G2_G2_G1_G1/FS_1/TEMP_P[0][1][0] ,
         \mat_kron/mult_40_G2_G2_G1_G1/A1[0] ,
         \mat_kron/mult_40_G2_G2_G1_G1/A1[1] ,
         \mat_kron/mult_40_G2_G2_G1_G1/A1[2] ,
         \mat_kron/mult_40_G2_G2_G1_G1/A1[3] ,
         \mat_kron/mult_40_G2_G2_G1_G1/A1[4] ,
         \mat_kron/mult_40_G2_G2_G1_G1/A1[5] ,
         \mat_kron/mult_40_G2_G2_G1_G1/A_notx[0] ,
         \mat_kron/mult_40_G2_G2_G1_G1/B_notx[0] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[0][1] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[0][2] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[0][3] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[0][4] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[0][5] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[0][6] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[0][7] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[1][0] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[1][1] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[1][2] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[1][3] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[1][4] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[1][5] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[1][6] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[2][0] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[2][1] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[2][2] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[2][3] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[2][4] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[2][5] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[3][0] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[3][1] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[3][2] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[3][3] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[3][4] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[4][0] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[4][1] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[4][2] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[4][3] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[5][0] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[5][1] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[5][2] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[6][0] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[6][1] ,
         \mat_kron/mult_40_G2_G2_G1_G1/ab[7][0] ,
         \mat_kron/mult_40_G2_G1/FS_1/P[0][0][1] ,
         \mat_kron/mult_40_G2_G1/FS_1/P[0][0][2] ,
         \mat_kron/mult_40_G2_G1/FS_1/P[0][0][3] ,
         \mat_kron/mult_40_G2_G1/FS_1/P[0][1][1] ,
         \mat_kron/mult_40_G2_G1/FS_1/TEMP_P[0][0][0] ,
         \mat_kron/mult_40_G2_G1/FS_1/TEMP_P[0][1][0] ,
         \mat_kron/mult_40_G2_G1/A1[0] , \mat_kron/mult_40_G2_G1/A1[1] ,
         \mat_kron/mult_40_G2_G1/A1[2] , \mat_kron/mult_40_G2_G1/A1[3] ,
         \mat_kron/mult_40_G2_G1/A1[4] , \mat_kron/mult_40_G2_G1/A1[5] ,
         \mat_kron/mult_40_G2_G1/A_notx[0] ,
         \mat_kron/mult_40_G2_G1/B_notx[0] , \mat_kron/mult_40_G2_G1/ab[0][1] ,
         \mat_kron/mult_40_G2_G1/ab[0][2] , \mat_kron/mult_40_G2_G1/ab[0][3] ,
         \mat_kron/mult_40_G2_G1/ab[0][4] , \mat_kron/mult_40_G2_G1/ab[0][5] ,
         \mat_kron/mult_40_G2_G1/ab[0][6] , \mat_kron/mult_40_G2_G1/ab[0][7] ,
         \mat_kron/mult_40_G2_G1/ab[1][0] , \mat_kron/mult_40_G2_G1/ab[1][1] ,
         \mat_kron/mult_40_G2_G1/ab[1][2] , \mat_kron/mult_40_G2_G1/ab[1][3] ,
         \mat_kron/mult_40_G2_G1/ab[1][4] , \mat_kron/mult_40_G2_G1/ab[1][5] ,
         \mat_kron/mult_40_G2_G1/ab[1][6] , \mat_kron/mult_40_G2_G1/ab[2][0] ,
         \mat_kron/mult_40_G2_G1/ab[2][1] , \mat_kron/mult_40_G2_G1/ab[2][2] ,
         \mat_kron/mult_40_G2_G1/ab[2][3] , \mat_kron/mult_40_G2_G1/ab[2][4] ,
         \mat_kron/mult_40_G2_G1/ab[2][5] , \mat_kron/mult_40_G2_G1/ab[3][0] ,
         \mat_kron/mult_40_G2_G1/ab[3][1] , \mat_kron/mult_40_G2_G1/ab[3][2] ,
         \mat_kron/mult_40_G2_G1/ab[3][3] , \mat_kron/mult_40_G2_G1/ab[3][4] ,
         \mat_kron/mult_40_G2_G1/ab[4][0] , \mat_kron/mult_40_G2_G1/ab[4][1] ,
         \mat_kron/mult_40_G2_G1/ab[4][2] , \mat_kron/mult_40_G2_G1/ab[4][3] ,
         \mat_kron/mult_40_G2_G1/ab[5][0] , \mat_kron/mult_40_G2_G1/ab[5][1] ,
         \mat_kron/mult_40_G2_G1/ab[5][2] , \mat_kron/mult_40_G2_G1/ab[6][0] ,
         \mat_kron/mult_40_G2_G1/ab[6][1] , \mat_kron/mult_40_G2_G1/ab[7][0] ,
         \mat_kron/mult_40_G2_G1_G2_G1/FS_1/P[0][0][1] ,
         \mat_kron/mult_40_G2_G1_G2_G1/FS_1/P[0][0][2] ,
         \mat_kron/mult_40_G2_G1_G2_G1/FS_1/P[0][0][3] ,
         \mat_kron/mult_40_G2_G1_G2_G1/FS_1/P[0][1][1] ,
         \mat_kron/mult_40_G2_G1_G2_G1/FS_1/TEMP_P[0][0][0] ,
         \mat_kron/mult_40_G2_G1_G2_G1/FS_1/TEMP_P[0][1][0] ,
         \mat_kron/mult_40_G2_G1_G2_G1/A1[0] ,
         \mat_kron/mult_40_G2_G1_G2_G1/A1[1] ,
         \mat_kron/mult_40_G2_G1_G2_G1/A1[2] ,
         \mat_kron/mult_40_G2_G1_G2_G1/A1[3] ,
         \mat_kron/mult_40_G2_G1_G2_G1/A1[4] ,
         \mat_kron/mult_40_G2_G1_G2_G1/A1[5] ,
         \mat_kron/mult_40_G2_G1_G2_G1/A_notx[0] ,
         \mat_kron/mult_40_G2_G1_G2_G1/B_notx[0] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[0][1] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[0][2] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[0][3] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[0][4] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[0][5] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[0][6] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[0][7] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[1][0] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[1][1] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[1][2] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[1][3] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[1][4] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[1][5] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[1][6] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[2][0] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[2][1] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[2][2] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[2][3] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[2][4] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[2][5] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[3][0] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[3][1] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[3][2] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[3][3] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[3][4] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[4][0] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[4][1] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[4][2] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[4][3] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[5][0] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[5][1] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[5][2] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[6][0] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[6][1] ,
         \mat_kron/mult_40_G2_G1_G2_G1/ab[7][0] ,
         \mat_kron/mult_40_G2_G2_G1/FS_1/P[0][0][1] ,
         \mat_kron/mult_40_G2_G2_G1/FS_1/P[0][0][2] ,
         \mat_kron/mult_40_G2_G2_G1/FS_1/P[0][0][3] ,
         \mat_kron/mult_40_G2_G2_G1/FS_1/P[0][1][1] ,
         \mat_kron/mult_40_G2_G2_G1/FS_1/TEMP_P[0][0][0] ,
         \mat_kron/mult_40_G2_G2_G1/FS_1/TEMP_P[0][1][0] ,
         \mat_kron/mult_40_G2_G2_G1/A1[0] , \mat_kron/mult_40_G2_G2_G1/A1[1] ,
         \mat_kron/mult_40_G2_G2_G1/A1[2] , \mat_kron/mult_40_G2_G2_G1/A1[3] ,
         \mat_kron/mult_40_G2_G2_G1/A1[4] , \mat_kron/mult_40_G2_G2_G1/A1[5] ,
         \mat_kron/mult_40_G2_G2_G1/A_notx[0] ,
         \mat_kron/mult_40_G2_G2_G1/B_notx[0] ,
         \mat_kron/mult_40_G2_G2_G1/ab[0][1] ,
         \mat_kron/mult_40_G2_G2_G1/ab[0][2] ,
         \mat_kron/mult_40_G2_G2_G1/ab[0][3] ,
         \mat_kron/mult_40_G2_G2_G1/ab[0][4] ,
         \mat_kron/mult_40_G2_G2_G1/ab[0][5] ,
         \mat_kron/mult_40_G2_G2_G1/ab[0][6] ,
         \mat_kron/mult_40_G2_G2_G1/ab[0][7] ,
         \mat_kron/mult_40_G2_G2_G1/ab[1][0] ,
         \mat_kron/mult_40_G2_G2_G1/ab[1][1] ,
         \mat_kron/mult_40_G2_G2_G1/ab[1][2] ,
         \mat_kron/mult_40_G2_G2_G1/ab[1][3] ,
         \mat_kron/mult_40_G2_G2_G1/ab[1][4] ,
         \mat_kron/mult_40_G2_G2_G1/ab[1][5] ,
         \mat_kron/mult_40_G2_G2_G1/ab[1][6] ,
         \mat_kron/mult_40_G2_G2_G1/ab[2][0] ,
         \mat_kron/mult_40_G2_G2_G1/ab[2][1] ,
         \mat_kron/mult_40_G2_G2_G1/ab[2][2] ,
         \mat_kron/mult_40_G2_G2_G1/ab[2][3] ,
         \mat_kron/mult_40_G2_G2_G1/ab[2][4] ,
         \mat_kron/mult_40_G2_G2_G1/ab[2][5] ,
         \mat_kron/mult_40_G2_G2_G1/ab[3][0] ,
         \mat_kron/mult_40_G2_G2_G1/ab[3][1] ,
         \mat_kron/mult_40_G2_G2_G1/ab[3][2] ,
         \mat_kron/mult_40_G2_G2_G1/ab[3][3] ,
         \mat_kron/mult_40_G2_G2_G1/ab[3][4] ,
         \mat_kron/mult_40_G2_G2_G1/ab[4][0] ,
         \mat_kron/mult_40_G2_G2_G1/ab[4][1] ,
         \mat_kron/mult_40_G2_G2_G1/ab[4][2] ,
         \mat_kron/mult_40_G2_G2_G1/ab[4][3] ,
         \mat_kron/mult_40_G2_G2_G1/ab[5][0] ,
         \mat_kron/mult_40_G2_G2_G1/ab[5][1] ,
         \mat_kron/mult_40_G2_G2_G1/ab[5][2] ,
         \mat_kron/mult_40_G2_G2_G1/ab[6][0] ,
         \mat_kron/mult_40_G2_G2_G1/ab[6][1] ,
         \mat_kron/mult_40_G2_G2_G1/ab[7][0] ,
         \mat_kron/mult_40_G2_G2_G2_G1/FS_1/P[0][0][1] ,
         \mat_kron/mult_40_G2_G2_G2_G1/FS_1/P[0][0][2] ,
         \mat_kron/mult_40_G2_G2_G2_G1/FS_1/P[0][0][3] ,
         \mat_kron/mult_40_G2_G2_G2_G1/FS_1/P[0][1][1] ,
         \mat_kron/mult_40_G2_G2_G2_G1/FS_1/TEMP_P[0][0][0] ,
         \mat_kron/mult_40_G2_G2_G2_G1/FS_1/TEMP_P[0][1][0] ,
         \mat_kron/mult_40_G2_G2_G2_G1/A1[0] ,
         \mat_kron/mult_40_G2_G2_G2_G1/A1[1] ,
         \mat_kron/mult_40_G2_G2_G2_G1/A1[2] ,
         \mat_kron/mult_40_G2_G2_G2_G1/A1[3] ,
         \mat_kron/mult_40_G2_G2_G2_G1/A1[4] ,
         \mat_kron/mult_40_G2_G2_G2_G1/A1[5] ,
         \mat_kron/mult_40_G2_G2_G2_G1/A_notx[0] ,
         \mat_kron/mult_40_G2_G2_G2_G1/B_notx[0] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[0][1] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[0][2] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[0][3] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[0][4] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[0][5] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[0][6] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[0][7] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[1][0] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[1][1] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[1][2] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[1][3] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[1][4] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[1][5] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[1][6] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[2][0] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[2][1] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[2][2] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[2][3] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[2][4] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[2][5] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[3][0] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[3][1] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[3][2] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[3][3] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[3][4] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[4][0] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[4][1] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[4][2] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[4][3] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[5][0] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[5][1] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[5][2] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[6][0] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[6][1] ,
         \mat_kron/mult_40_G2_G2_G2_G1/ab[7][0] ,
         \mat_kron/mult_40_G2/FS_1/P[0][0][1] ,
         \mat_kron/mult_40_G2/FS_1/P[0][0][2] ,
         \mat_kron/mult_40_G2/FS_1/P[0][0][3] ,
         \mat_kron/mult_40_G2/FS_1/P[0][1][1] ,
         \mat_kron/mult_40_G2/FS_1/TEMP_P[0][0][0] ,
         \mat_kron/mult_40_G2/FS_1/TEMP_P[0][1][0] ,
         \mat_kron/mult_40_G2/A1[0] , \mat_kron/mult_40_G2/A1[1] ,
         \mat_kron/mult_40_G2/A1[2] , \mat_kron/mult_40_G2/A1[3] ,
         \mat_kron/mult_40_G2/A1[4] , \mat_kron/mult_40_G2/A1[5] ,
         \mat_kron/mult_40_G2/A_notx[0] , \mat_kron/mult_40_G2/B_notx[0] ,
         \mat_kron/mult_40_G2/ab[0][1] , \mat_kron/mult_40_G2/ab[0][2] ,
         \mat_kron/mult_40_G2/ab[0][3] , \mat_kron/mult_40_G2/ab[0][4] ,
         \mat_kron/mult_40_G2/ab[0][5] , \mat_kron/mult_40_G2/ab[0][6] ,
         \mat_kron/mult_40_G2/ab[0][7] , \mat_kron/mult_40_G2/ab[1][0] ,
         \mat_kron/mult_40_G2/ab[1][1] , \mat_kron/mult_40_G2/ab[1][2] ,
         \mat_kron/mult_40_G2/ab[1][3] , \mat_kron/mult_40_G2/ab[1][4] ,
         \mat_kron/mult_40_G2/ab[1][5] , \mat_kron/mult_40_G2/ab[1][6] ,
         \mat_kron/mult_40_G2/ab[2][0] , \mat_kron/mult_40_G2/ab[2][1] ,
         \mat_kron/mult_40_G2/ab[2][2] , \mat_kron/mult_40_G2/ab[2][3] ,
         \mat_kron/mult_40_G2/ab[2][4] , \mat_kron/mult_40_G2/ab[2][5] ,
         \mat_kron/mult_40_G2/ab[3][0] , \mat_kron/mult_40_G2/ab[3][1] ,
         \mat_kron/mult_40_G2/ab[3][2] , \mat_kron/mult_40_G2/ab[3][3] ,
         \mat_kron/mult_40_G2/ab[3][4] , \mat_kron/mult_40_G2/ab[4][0] ,
         \mat_kron/mult_40_G2/ab[4][1] , \mat_kron/mult_40_G2/ab[4][2] ,
         \mat_kron/mult_40_G2/ab[4][3] , \mat_kron/mult_40_G2/ab[5][0] ,
         \mat_kron/mult_40_G2/ab[5][1] , \mat_kron/mult_40_G2/ab[5][2] ,
         \mat_kron/mult_40_G2/ab[6][0] , \mat_kron/mult_40_G2/ab[6][1] ,
         \mat_kron/mult_40_G2/ab[7][0] ,
         \mat_kron/mult_40_G2_G1_G1_G2/FS_1/P[0][0][1] ,
         \mat_kron/mult_40_G2_G1_G1_G2/FS_1/P[0][0][2] ,
         \mat_kron/mult_40_G2_G1_G1_G2/FS_1/P[0][0][3] ,
         \mat_kron/mult_40_G2_G1_G1_G2/FS_1/P[0][1][1] ,
         \mat_kron/mult_40_G2_G1_G1_G2/FS_1/TEMP_P[0][0][0] ,
         \mat_kron/mult_40_G2_G1_G1_G2/FS_1/TEMP_P[0][1][0] ,
         \mat_kron/mult_40_G2_G1_G1_G2/A1[0] ,
         \mat_kron/mult_40_G2_G1_G1_G2/A1[1] ,
         \mat_kron/mult_40_G2_G1_G1_G2/A1[2] ,
         \mat_kron/mult_40_G2_G1_G1_G2/A1[3] ,
         \mat_kron/mult_40_G2_G1_G1_G2/A1[4] ,
         \mat_kron/mult_40_G2_G1_G1_G2/A1[5] ,
         \mat_kron/mult_40_G2_G1_G1_G2/A_notx[0] ,
         \mat_kron/mult_40_G2_G1_G1_G2/B_notx[0] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[0][1] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[0][2] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[0][3] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[0][4] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[0][5] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[0][6] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[0][7] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[1][0] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[1][1] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[1][2] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[1][3] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[1][4] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[1][5] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[1][6] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[2][0] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[2][1] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[2][2] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[2][3] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[2][4] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[2][5] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[3][0] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[3][1] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[3][2] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[3][3] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[3][4] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[4][0] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[4][1] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[4][2] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[4][3] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[5][0] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[5][1] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[5][2] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[6][0] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[6][1] ,
         \mat_kron/mult_40_G2_G1_G1_G2/ab[7][0] ,
         \mat_kron/mult_40_G2_G1_G2/FS_1/P[0][0][1] ,
         \mat_kron/mult_40_G2_G1_G2/FS_1/P[0][0][2] ,
         \mat_kron/mult_40_G2_G1_G2/FS_1/P[0][0][3] ,
         \mat_kron/mult_40_G2_G1_G2/FS_1/P[0][1][1] ,
         \mat_kron/mult_40_G2_G1_G2/FS_1/TEMP_P[0][0][0] ,
         \mat_kron/mult_40_G2_G1_G2/FS_1/TEMP_P[0][1][0] ,
         \mat_kron/mult_40_G2_G1_G2/A1[0] , \mat_kron/mult_40_G2_G1_G2/A1[1] ,
         \mat_kron/mult_40_G2_G1_G2/A1[2] , \mat_kron/mult_40_G2_G1_G2/A1[3] ,
         \mat_kron/mult_40_G2_G1_G2/A1[4] , \mat_kron/mult_40_G2_G1_G2/A1[5] ,
         \mat_kron/mult_40_G2_G1_G2/A_notx[0] ,
         \mat_kron/mult_40_G2_G1_G2/B_notx[0] ,
         \mat_kron/mult_40_G2_G1_G2/ab[0][1] ,
         \mat_kron/mult_40_G2_G1_G2/ab[0][2] ,
         \mat_kron/mult_40_G2_G1_G2/ab[0][3] ,
         \mat_kron/mult_40_G2_G1_G2/ab[0][4] ,
         \mat_kron/mult_40_G2_G1_G2/ab[0][5] ,
         \mat_kron/mult_40_G2_G1_G2/ab[0][6] ,
         \mat_kron/mult_40_G2_G1_G2/ab[0][7] ,
         \mat_kron/mult_40_G2_G1_G2/ab[1][0] ,
         \mat_kron/mult_40_G2_G1_G2/ab[1][1] ,
         \mat_kron/mult_40_G2_G1_G2/ab[1][2] ,
         \mat_kron/mult_40_G2_G1_G2/ab[1][3] ,
         \mat_kron/mult_40_G2_G1_G2/ab[1][4] ,
         \mat_kron/mult_40_G2_G1_G2/ab[1][5] ,
         \mat_kron/mult_40_G2_G1_G2/ab[1][6] ,
         \mat_kron/mult_40_G2_G1_G2/ab[2][0] ,
         \mat_kron/mult_40_G2_G1_G2/ab[2][1] ,
         \mat_kron/mult_40_G2_G1_G2/ab[2][2] ,
         \mat_kron/mult_40_G2_G1_G2/ab[2][3] ,
         \mat_kron/mult_40_G2_G1_G2/ab[2][4] ,
         \mat_kron/mult_40_G2_G1_G2/ab[2][5] ,
         \mat_kron/mult_40_G2_G1_G2/ab[3][0] ,
         \mat_kron/mult_40_G2_G1_G2/ab[3][1] ,
         \mat_kron/mult_40_G2_G1_G2/ab[3][2] ,
         \mat_kron/mult_40_G2_G1_G2/ab[3][3] ,
         \mat_kron/mult_40_G2_G1_G2/ab[3][4] ,
         \mat_kron/mult_40_G2_G1_G2/ab[4][0] ,
         \mat_kron/mult_40_G2_G1_G2/ab[4][1] ,
         \mat_kron/mult_40_G2_G1_G2/ab[4][2] ,
         \mat_kron/mult_40_G2_G1_G2/ab[4][3] ,
         \mat_kron/mult_40_G2_G1_G2/ab[5][0] ,
         \mat_kron/mult_40_G2_G1_G2/ab[5][1] ,
         \mat_kron/mult_40_G2_G1_G2/ab[5][2] ,
         \mat_kron/mult_40_G2_G1_G2/ab[6][0] ,
         \mat_kron/mult_40_G2_G1_G2/ab[6][1] ,
         \mat_kron/mult_40_G2_G1_G2/ab[7][0] ,
         \mat_kron/mult_40_G2_G2_G1_G2/FS_1/P[0][0][1] ,
         \mat_kron/mult_40_G2_G2_G1_G2/FS_1/P[0][0][2] ,
         \mat_kron/mult_40_G2_G2_G1_G2/FS_1/P[0][0][3] ,
         \mat_kron/mult_40_G2_G2_G1_G2/FS_1/P[0][1][1] ,
         \mat_kron/mult_40_G2_G2_G1_G2/FS_1/TEMP_P[0][0][0] ,
         \mat_kron/mult_40_G2_G2_G1_G2/FS_1/TEMP_P[0][1][0] ,
         \mat_kron/mult_40_G2_G2_G1_G2/A1[0] ,
         \mat_kron/mult_40_G2_G2_G1_G2/A1[1] ,
         \mat_kron/mult_40_G2_G2_G1_G2/A1[2] ,
         \mat_kron/mult_40_G2_G2_G1_G2/A1[3] ,
         \mat_kron/mult_40_G2_G2_G1_G2/A1[4] ,
         \mat_kron/mult_40_G2_G2_G1_G2/A1[5] ,
         \mat_kron/mult_40_G2_G2_G1_G2/A_notx[0] ,
         \mat_kron/mult_40_G2_G2_G1_G2/B_notx[0] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[0][1] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[0][2] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[0][3] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[0][4] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[0][5] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[0][6] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[0][7] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[1][0] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[1][1] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[1][2] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[1][3] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[1][4] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[1][5] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[1][6] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[2][0] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[2][1] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[2][2] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[2][3] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[2][4] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[2][5] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[3][0] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[3][1] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[3][2] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[3][3] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[3][4] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[4][0] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[4][1] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[4][2] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[4][3] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[5][0] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[5][1] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[5][2] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[6][0] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[6][1] ,
         \mat_kron/mult_40_G2_G2_G1_G2/ab[7][0] ,
         \mat_kron/mult_40_G2_G2/FS_1/P[0][0][1] ,
         \mat_kron/mult_40_G2_G2/FS_1/P[0][0][2] ,
         \mat_kron/mult_40_G2_G2/FS_1/P[0][0][3] ,
         \mat_kron/mult_40_G2_G2/FS_1/P[0][1][1] ,
         \mat_kron/mult_40_G2_G2/FS_1/TEMP_P[0][0][0] ,
         \mat_kron/mult_40_G2_G2/FS_1/TEMP_P[0][1][0] ,
         \mat_kron/mult_40_G2_G2/A1[0] , \mat_kron/mult_40_G2_G2/A1[1] ,
         \mat_kron/mult_40_G2_G2/A1[2] , \mat_kron/mult_40_G2_G2/A1[3] ,
         \mat_kron/mult_40_G2_G2/A1[4] , \mat_kron/mult_40_G2_G2/A1[5] ,
         \mat_kron/mult_40_G2_G2/A_notx[0] ,
         \mat_kron/mult_40_G2_G2/B_notx[0] , \mat_kron/mult_40_G2_G2/ab[0][1] ,
         \mat_kron/mult_40_G2_G2/ab[0][2] , \mat_kron/mult_40_G2_G2/ab[0][3] ,
         \mat_kron/mult_40_G2_G2/ab[0][4] , \mat_kron/mult_40_G2_G2/ab[0][5] ,
         \mat_kron/mult_40_G2_G2/ab[0][6] , \mat_kron/mult_40_G2_G2/ab[0][7] ,
         \mat_kron/mult_40_G2_G2/ab[1][0] , \mat_kron/mult_40_G2_G2/ab[1][1] ,
         \mat_kron/mult_40_G2_G2/ab[1][2] , \mat_kron/mult_40_G2_G2/ab[1][3] ,
         \mat_kron/mult_40_G2_G2/ab[1][4] , \mat_kron/mult_40_G2_G2/ab[1][5] ,
         \mat_kron/mult_40_G2_G2/ab[1][6] , \mat_kron/mult_40_G2_G2/ab[2][0] ,
         \mat_kron/mult_40_G2_G2/ab[2][1] , \mat_kron/mult_40_G2_G2/ab[2][2] ,
         \mat_kron/mult_40_G2_G2/ab[2][3] , \mat_kron/mult_40_G2_G2/ab[2][4] ,
         \mat_kron/mult_40_G2_G2/ab[2][5] , \mat_kron/mult_40_G2_G2/ab[3][0] ,
         \mat_kron/mult_40_G2_G2/ab[3][1] , \mat_kron/mult_40_G2_G2/ab[3][2] ,
         \mat_kron/mult_40_G2_G2/ab[3][3] , \mat_kron/mult_40_G2_G2/ab[3][4] ,
         \mat_kron/mult_40_G2_G2/ab[4][0] , \mat_kron/mult_40_G2_G2/ab[4][1] ,
         \mat_kron/mult_40_G2_G2/ab[4][2] , \mat_kron/mult_40_G2_G2/ab[4][3] ,
         \mat_kron/mult_40_G2_G2/ab[5][0] , \mat_kron/mult_40_G2_G2/ab[5][1] ,
         \mat_kron/mult_40_G2_G2/ab[5][2] , \mat_kron/mult_40_G2_G2/ab[6][0] ,
         \mat_kron/mult_40_G2_G2/ab[6][1] , \mat_kron/mult_40_G2_G2/ab[7][0] ,
         \mat_kron/mult_40_G2_G1_G2_G2/FS_1/P[0][0][1] ,
         \mat_kron/mult_40_G2_G1_G2_G2/FS_1/P[0][0][2] ,
         \mat_kron/mult_40_G2_G1_G2_G2/FS_1/P[0][0][3] ,
         \mat_kron/mult_40_G2_G1_G2_G2/FS_1/P[0][1][1] ,
         \mat_kron/mult_40_G2_G1_G2_G2/FS_1/TEMP_P[0][0][0] ,
         \mat_kron/mult_40_G2_G1_G2_G2/FS_1/TEMP_P[0][1][0] ,
         \mat_kron/mult_40_G2_G1_G2_G2/A1[0] ,
         \mat_kron/mult_40_G2_G1_G2_G2/A1[1] ,
         \mat_kron/mult_40_G2_G1_G2_G2/A1[2] ,
         \mat_kron/mult_40_G2_G1_G2_G2/A1[3] ,
         \mat_kron/mult_40_G2_G1_G2_G2/A1[4] ,
         \mat_kron/mult_40_G2_G1_G2_G2/A1[5] ,
         \mat_kron/mult_40_G2_G1_G2_G2/A_notx[0] ,
         \mat_kron/mult_40_G2_G1_G2_G2/B_notx[0] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[0][1] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[0][2] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[0][3] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[0][4] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[0][5] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[0][6] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[0][7] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[1][0] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[1][1] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[1][2] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[1][3] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[1][4] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[1][5] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[1][6] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[2][0] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[2][1] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[2][2] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[2][3] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[2][4] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[2][5] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[3][0] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[3][1] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[3][2] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[3][3] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[3][4] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[4][0] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[4][1] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[4][2] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[4][3] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[5][0] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[5][1] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[5][2] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[6][0] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[6][1] ,
         \mat_kron/mult_40_G2_G1_G2_G2/ab[7][0] ,
         \mat_kron/mult_40_G2_G2_G2/FS_1/P[0][0][1] ,
         \mat_kron/mult_40_G2_G2_G2/FS_1/P[0][0][2] ,
         \mat_kron/mult_40_G2_G2_G2/FS_1/P[0][0][3] ,
         \mat_kron/mult_40_G2_G2_G2/FS_1/P[0][1][1] ,
         \mat_kron/mult_40_G2_G2_G2/FS_1/TEMP_P[0][0][0] ,
         \mat_kron/mult_40_G2_G2_G2/FS_1/TEMP_P[0][1][0] ,
         \mat_kron/mult_40_G2_G2_G2/A1[0] , \mat_kron/mult_40_G2_G2_G2/A1[1] ,
         \mat_kron/mult_40_G2_G2_G2/A1[2] , \mat_kron/mult_40_G2_G2_G2/A1[3] ,
         \mat_kron/mult_40_G2_G2_G2/A1[4] , \mat_kron/mult_40_G2_G2_G2/A1[5] ,
         \mat_kron/mult_40_G2_G2_G2/A_notx[0] ,
         \mat_kron/mult_40_G2_G2_G2/B_notx[0] ,
         \mat_kron/mult_40_G2_G2_G2/ab[0][1] ,
         \mat_kron/mult_40_G2_G2_G2/ab[0][2] ,
         \mat_kron/mult_40_G2_G2_G2/ab[0][3] ,
         \mat_kron/mult_40_G2_G2_G2/ab[0][4] ,
         \mat_kron/mult_40_G2_G2_G2/ab[0][5] ,
         \mat_kron/mult_40_G2_G2_G2/ab[0][6] ,
         \mat_kron/mult_40_G2_G2_G2/ab[0][7] ,
         \mat_kron/mult_40_G2_G2_G2/ab[1][0] ,
         \mat_kron/mult_40_G2_G2_G2/ab[1][1] ,
         \mat_kron/mult_40_G2_G2_G2/ab[1][2] ,
         \mat_kron/mult_40_G2_G2_G2/ab[1][3] ,
         \mat_kron/mult_40_G2_G2_G2/ab[1][4] ,
         \mat_kron/mult_40_G2_G2_G2/ab[1][5] ,
         \mat_kron/mult_40_G2_G2_G2/ab[1][6] ,
         \mat_kron/mult_40_G2_G2_G2/ab[2][0] ,
         \mat_kron/mult_40_G2_G2_G2/ab[2][1] ,
         \mat_kron/mult_40_G2_G2_G2/ab[2][2] ,
         \mat_kron/mult_40_G2_G2_G2/ab[2][3] ,
         \mat_kron/mult_40_G2_G2_G2/ab[2][4] ,
         \mat_kron/mult_40_G2_G2_G2/ab[2][5] ,
         \mat_kron/mult_40_G2_G2_G2/ab[3][0] ,
         \mat_kron/mult_40_G2_G2_G2/ab[3][1] ,
         \mat_kron/mult_40_G2_G2_G2/ab[3][2] ,
         \mat_kron/mult_40_G2_G2_G2/ab[3][3] ,
         \mat_kron/mult_40_G2_G2_G2/ab[3][4] ,
         \mat_kron/mult_40_G2_G2_G2/ab[4][0] ,
         \mat_kron/mult_40_G2_G2_G2/ab[4][1] ,
         \mat_kron/mult_40_G2_G2_G2/ab[4][2] ,
         \mat_kron/mult_40_G2_G2_G2/ab[4][3] ,
         \mat_kron/mult_40_G2_G2_G2/ab[5][0] ,
         \mat_kron/mult_40_G2_G2_G2/ab[5][1] ,
         \mat_kron/mult_40_G2_G2_G2/ab[5][2] ,
         \mat_kron/mult_40_G2_G2_G2/ab[6][0] ,
         \mat_kron/mult_40_G2_G2_G2/ab[6][1] ,
         \mat_kron/mult_40_G2_G2_G2/ab[7][0] ,
         \mat_kron/mult_40_G2_G2_G2_G2/FS_1/P[0][0][1] ,
         \mat_kron/mult_40_G2_G2_G2_G2/FS_1/P[0][0][2] ,
         \mat_kron/mult_40_G2_G2_G2_G2/FS_1/P[0][0][3] ,
         \mat_kron/mult_40_G2_G2_G2_G2/FS_1/P[0][1][1] ,
         \mat_kron/mult_40_G2_G2_G2_G2/FS_1/TEMP_P[0][0][0] ,
         \mat_kron/mult_40_G2_G2_G2_G2/FS_1/TEMP_P[0][1][0] ,
         \mat_kron/mult_40_G2_G2_G2_G2/A1[0] ,
         \mat_kron/mult_40_G2_G2_G2_G2/A1[1] ,
         \mat_kron/mult_40_G2_G2_G2_G2/A1[2] ,
         \mat_kron/mult_40_G2_G2_G2_G2/A1[3] ,
         \mat_kron/mult_40_G2_G2_G2_G2/A1[4] ,
         \mat_kron/mult_40_G2_G2_G2_G2/A1[5] ,
         \mat_kron/mult_40_G2_G2_G2_G2/A_notx[0] ,
         \mat_kron/mult_40_G2_G2_G2_G2/B_notx[0] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[0][1] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[0][2] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[0][3] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[0][4] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[0][5] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[0][6] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[0][7] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[1][0] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[1][1] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[1][2] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[1][3] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[1][4] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[1][5] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[1][6] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[2][0] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[2][1] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[2][2] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[2][3] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[2][4] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[2][5] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[3][0] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[3][1] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[3][2] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[3][3] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[3][4] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[4][0] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[4][1] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[4][2] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[4][3] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[5][0] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[5][1] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[5][2] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[6][0] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[6][1] ,
         \mat_kron/mult_40_G2_G2_G2_G2/ab[7][0] ,
         \mat_mul/mult_37/FS_1/P[0][0][1] , \mat_mul/mult_37/FS_1/P[0][0][2] ,
         \mat_mul/mult_37/FS_1/P[0][0][3] , \mat_mul/mult_37/FS_1/P[0][1][1] ,
         \mat_mul/mult_37/FS_1/TEMP_P[0][0][0] ,
         \mat_mul/mult_37/FS_1/TEMP_P[0][1][0] , \mat_mul/mult_37/A1[0] ,
         \mat_mul/mult_37/A1[1] , \mat_mul/mult_37/A1[2] ,
         \mat_mul/mult_37/A1[3] , \mat_mul/mult_37/A1[4] ,
         \mat_mul/mult_37/A1[5] , \mat_mul/mult_37/A_notx[0] ,
         \mat_mul/mult_37/B_notx[0] , \mat_mul/mult_37/ab[0][1] ,
         \mat_mul/mult_37/ab[0][2] , \mat_mul/mult_37/ab[0][3] ,
         \mat_mul/mult_37/ab[0][4] , \mat_mul/mult_37/ab[0][5] ,
         \mat_mul/mult_37/ab[0][6] , \mat_mul/mult_37/ab[0][7] ,
         \mat_mul/mult_37/ab[1][0] , \mat_mul/mult_37/ab[1][1] ,
         \mat_mul/mult_37/ab[1][2] , \mat_mul/mult_37/ab[1][3] ,
         \mat_mul/mult_37/ab[1][4] , \mat_mul/mult_37/ab[1][5] ,
         \mat_mul/mult_37/ab[1][6] , \mat_mul/mult_37/ab[2][0] ,
         \mat_mul/mult_37/ab[2][1] , \mat_mul/mult_37/ab[2][2] ,
         \mat_mul/mult_37/ab[2][3] , \mat_mul/mult_37/ab[2][4] ,
         \mat_mul/mult_37/ab[2][5] , \mat_mul/mult_37/ab[3][0] ,
         \mat_mul/mult_37/ab[3][1] , \mat_mul/mult_37/ab[3][2] ,
         \mat_mul/mult_37/ab[3][3] , \mat_mul/mult_37/ab[3][4] ,
         \mat_mul/mult_37/ab[4][0] , \mat_mul/mult_37/ab[4][1] ,
         \mat_mul/mult_37/ab[4][2] , \mat_mul/mult_37/ab[4][3] ,
         \mat_mul/mult_37/ab[5][0] , \mat_mul/mult_37/ab[5][1] ,
         \mat_mul/mult_37/ab[5][2] , \mat_mul/mult_37/ab[6][0] ,
         \mat_mul/mult_37/ab[6][1] , \mat_mul/mult_37/ab[7][0] ,
         \mat_mul/mult_37_G2_G1_G1/FS_1/P[0][0][1] ,
         \mat_mul/mult_37_G2_G1_G1/FS_1/P[0][0][2] ,
         \mat_mul/mult_37_G2_G1_G1/FS_1/P[0][0][3] ,
         \mat_mul/mult_37_G2_G1_G1/FS_1/P[0][1][1] ,
         \mat_mul/mult_37_G2_G1_G1/FS_1/TEMP_P[0][0][0] ,
         \mat_mul/mult_37_G2_G1_G1/FS_1/TEMP_P[0][1][0] ,
         \mat_mul/mult_37_G2_G1_G1/A1[0] , \mat_mul/mult_37_G2_G1_G1/A1[1] ,
         \mat_mul/mult_37_G2_G1_G1/A1[2] , \mat_mul/mult_37_G2_G1_G1/A1[3] ,
         \mat_mul/mult_37_G2_G1_G1/A1[4] , \mat_mul/mult_37_G2_G1_G1/A1[5] ,
         \mat_mul/mult_37_G2_G1_G1/A_notx[0] ,
         \mat_mul/mult_37_G2_G1_G1/B_notx[0] ,
         \mat_mul/mult_37_G2_G1_G1/ab[0][1] ,
         \mat_mul/mult_37_G2_G1_G1/ab[0][2] ,
         \mat_mul/mult_37_G2_G1_G1/ab[0][3] ,
         \mat_mul/mult_37_G2_G1_G1/ab[0][4] ,
         \mat_mul/mult_37_G2_G1_G1/ab[0][5] ,
         \mat_mul/mult_37_G2_G1_G1/ab[0][6] ,
         \mat_mul/mult_37_G2_G1_G1/ab[0][7] ,
         \mat_mul/mult_37_G2_G1_G1/ab[1][0] ,
         \mat_mul/mult_37_G2_G1_G1/ab[1][1] ,
         \mat_mul/mult_37_G2_G1_G1/ab[1][2] ,
         \mat_mul/mult_37_G2_G1_G1/ab[1][3] ,
         \mat_mul/mult_37_G2_G1_G1/ab[1][4] ,
         \mat_mul/mult_37_G2_G1_G1/ab[1][5] ,
         \mat_mul/mult_37_G2_G1_G1/ab[1][6] ,
         \mat_mul/mult_37_G2_G1_G1/ab[2][0] ,
         \mat_mul/mult_37_G2_G1_G1/ab[2][1] ,
         \mat_mul/mult_37_G2_G1_G1/ab[2][2] ,
         \mat_mul/mult_37_G2_G1_G1/ab[2][3] ,
         \mat_mul/mult_37_G2_G1_G1/ab[2][4] ,
         \mat_mul/mult_37_G2_G1_G1/ab[2][5] ,
         \mat_mul/mult_37_G2_G1_G1/ab[3][0] ,
         \mat_mul/mult_37_G2_G1_G1/ab[3][1] ,
         \mat_mul/mult_37_G2_G1_G1/ab[3][2] ,
         \mat_mul/mult_37_G2_G1_G1/ab[3][3] ,
         \mat_mul/mult_37_G2_G1_G1/ab[3][4] ,
         \mat_mul/mult_37_G2_G1_G1/ab[4][0] ,
         \mat_mul/mult_37_G2_G1_G1/ab[4][1] ,
         \mat_mul/mult_37_G2_G1_G1/ab[4][2] ,
         \mat_mul/mult_37_G2_G1_G1/ab[4][3] ,
         \mat_mul/mult_37_G2_G1_G1/ab[5][0] ,
         \mat_mul/mult_37_G2_G1_G1/ab[5][1] ,
         \mat_mul/mult_37_G2_G1_G1/ab[5][2] ,
         \mat_mul/mult_37_G2_G1_G1/ab[6][0] ,
         \mat_mul/mult_37_G2_G1_G1/ab[6][1] ,
         \mat_mul/mult_37_G2_G1_G1/ab[7][0] ,
         \mat_mul/mult_37_G2_G1/FS_1/P[0][0][1] ,
         \mat_mul/mult_37_G2_G1/FS_1/P[0][0][2] ,
         \mat_mul/mult_37_G2_G1/FS_1/P[0][0][3] ,
         \mat_mul/mult_37_G2_G1/FS_1/P[0][1][1] ,
         \mat_mul/mult_37_G2_G1/FS_1/TEMP_P[0][0][0] ,
         \mat_mul/mult_37_G2_G1/FS_1/TEMP_P[0][1][0] ,
         \mat_mul/mult_37_G2_G1/A1[0] , \mat_mul/mult_37_G2_G1/A1[1] ,
         \mat_mul/mult_37_G2_G1/A1[2] , \mat_mul/mult_37_G2_G1/A1[3] ,
         \mat_mul/mult_37_G2_G1/A1[4] , \mat_mul/mult_37_G2_G1/A1[5] ,
         \mat_mul/mult_37_G2_G1/A_notx[0] , \mat_mul/mult_37_G2_G1/B_notx[0] ,
         \mat_mul/mult_37_G2_G1/ab[0][1] , \mat_mul/mult_37_G2_G1/ab[0][2] ,
         \mat_mul/mult_37_G2_G1/ab[0][3] , \mat_mul/mult_37_G2_G1/ab[0][4] ,
         \mat_mul/mult_37_G2_G1/ab[0][5] , \mat_mul/mult_37_G2_G1/ab[0][6] ,
         \mat_mul/mult_37_G2_G1/ab[0][7] , \mat_mul/mult_37_G2_G1/ab[1][0] ,
         \mat_mul/mult_37_G2_G1/ab[1][1] , \mat_mul/mult_37_G2_G1/ab[1][2] ,
         \mat_mul/mult_37_G2_G1/ab[1][3] , \mat_mul/mult_37_G2_G1/ab[1][4] ,
         \mat_mul/mult_37_G2_G1/ab[1][5] , \mat_mul/mult_37_G2_G1/ab[1][6] ,
         \mat_mul/mult_37_G2_G1/ab[2][0] , \mat_mul/mult_37_G2_G1/ab[2][1] ,
         \mat_mul/mult_37_G2_G1/ab[2][2] , \mat_mul/mult_37_G2_G1/ab[2][3] ,
         \mat_mul/mult_37_G2_G1/ab[2][4] , \mat_mul/mult_37_G2_G1/ab[2][5] ,
         \mat_mul/mult_37_G2_G1/ab[3][0] , \mat_mul/mult_37_G2_G1/ab[3][1] ,
         \mat_mul/mult_37_G2_G1/ab[3][2] , \mat_mul/mult_37_G2_G1/ab[3][3] ,
         \mat_mul/mult_37_G2_G1/ab[3][4] , \mat_mul/mult_37_G2_G1/ab[4][0] ,
         \mat_mul/mult_37_G2_G1/ab[4][1] , \mat_mul/mult_37_G2_G1/ab[4][2] ,
         \mat_mul/mult_37_G2_G1/ab[4][3] , \mat_mul/mult_37_G2_G1/ab[5][0] ,
         \mat_mul/mult_37_G2_G1/ab[5][1] , \mat_mul/mult_37_G2_G1/ab[5][2] ,
         \mat_mul/mult_37_G2_G1/ab[6][0] , \mat_mul/mult_37_G2_G1/ab[6][1] ,
         \mat_mul/mult_37_G2_G1/ab[7][0] ,
         \mat_mul/mult_37_G2_G2_G1/FS_1/P[0][0][1] ,
         \mat_mul/mult_37_G2_G2_G1/FS_1/P[0][0][2] ,
         \mat_mul/mult_37_G2_G2_G1/FS_1/P[0][0][3] ,
         \mat_mul/mult_37_G2_G2_G1/FS_1/P[0][1][1] ,
         \mat_mul/mult_37_G2_G2_G1/FS_1/TEMP_P[0][0][0] ,
         \mat_mul/mult_37_G2_G2_G1/FS_1/TEMP_P[0][1][0] ,
         \mat_mul/mult_37_G2_G2_G1/A1[0] , \mat_mul/mult_37_G2_G2_G1/A1[1] ,
         \mat_mul/mult_37_G2_G2_G1/A1[2] , \mat_mul/mult_37_G2_G2_G1/A1[3] ,
         \mat_mul/mult_37_G2_G2_G1/A1[4] , \mat_mul/mult_37_G2_G2_G1/A1[5] ,
         \mat_mul/mult_37_G2_G2_G1/A_notx[0] ,
         \mat_mul/mult_37_G2_G2_G1/B_notx[0] ,
         \mat_mul/mult_37_G2_G2_G1/ab[0][1] ,
         \mat_mul/mult_37_G2_G2_G1/ab[0][2] ,
         \mat_mul/mult_37_G2_G2_G1/ab[0][3] ,
         \mat_mul/mult_37_G2_G2_G1/ab[0][4] ,
         \mat_mul/mult_37_G2_G2_G1/ab[0][5] ,
         \mat_mul/mult_37_G2_G2_G1/ab[0][6] ,
         \mat_mul/mult_37_G2_G2_G1/ab[0][7] ,
         \mat_mul/mult_37_G2_G2_G1/ab[1][0] ,
         \mat_mul/mult_37_G2_G2_G1/ab[1][1] ,
         \mat_mul/mult_37_G2_G2_G1/ab[1][2] ,
         \mat_mul/mult_37_G2_G2_G1/ab[1][3] ,
         \mat_mul/mult_37_G2_G2_G1/ab[1][4] ,
         \mat_mul/mult_37_G2_G2_G1/ab[1][5] ,
         \mat_mul/mult_37_G2_G2_G1/ab[1][6] ,
         \mat_mul/mult_37_G2_G2_G1/ab[2][0] ,
         \mat_mul/mult_37_G2_G2_G1/ab[2][1] ,
         \mat_mul/mult_37_G2_G2_G1/ab[2][2] ,
         \mat_mul/mult_37_G2_G2_G1/ab[2][3] ,
         \mat_mul/mult_37_G2_G2_G1/ab[2][4] ,
         \mat_mul/mult_37_G2_G2_G1/ab[2][5] ,
         \mat_mul/mult_37_G2_G2_G1/ab[3][0] ,
         \mat_mul/mult_37_G2_G2_G1/ab[3][1] ,
         \mat_mul/mult_37_G2_G2_G1/ab[3][2] ,
         \mat_mul/mult_37_G2_G2_G1/ab[3][3] ,
         \mat_mul/mult_37_G2_G2_G1/ab[3][4] ,
         \mat_mul/mult_37_G2_G2_G1/ab[4][0] ,
         \mat_mul/mult_37_G2_G2_G1/ab[4][1] ,
         \mat_mul/mult_37_G2_G2_G1/ab[4][2] ,
         \mat_mul/mult_37_G2_G2_G1/ab[4][3] ,
         \mat_mul/mult_37_G2_G2_G1/ab[5][0] ,
         \mat_mul/mult_37_G2_G2_G1/ab[5][1] ,
         \mat_mul/mult_37_G2_G2_G1/ab[5][2] ,
         \mat_mul/mult_37_G2_G2_G1/ab[6][0] ,
         \mat_mul/mult_37_G2_G2_G1/ab[6][1] ,
         \mat_mul/mult_37_G2_G2_G1/ab[7][0] ,
         \mat_mul/mult_37_G2/FS_1/P[0][0][1] ,
         \mat_mul/mult_37_G2/FS_1/P[0][0][2] ,
         \mat_mul/mult_37_G2/FS_1/P[0][0][3] ,
         \mat_mul/mult_37_G2/FS_1/P[0][1][1] ,
         \mat_mul/mult_37_G2/FS_1/TEMP_P[0][0][0] ,
         \mat_mul/mult_37_G2/FS_1/TEMP_P[0][1][0] , \mat_mul/mult_37_G2/A1[0] ,
         \mat_mul/mult_37_G2/A1[1] , \mat_mul/mult_37_G2/A1[2] ,
         \mat_mul/mult_37_G2/A1[3] , \mat_mul/mult_37_G2/A1[4] ,
         \mat_mul/mult_37_G2/A1[5] , \mat_mul/mult_37_G2/A_notx[0] ,
         \mat_mul/mult_37_G2/B_notx[0] , \mat_mul/mult_37_G2/ab[0][1] ,
         \mat_mul/mult_37_G2/ab[0][2] , \mat_mul/mult_37_G2/ab[0][3] ,
         \mat_mul/mult_37_G2/ab[0][4] , \mat_mul/mult_37_G2/ab[0][5] ,
         \mat_mul/mult_37_G2/ab[0][6] , \mat_mul/mult_37_G2/ab[0][7] ,
         \mat_mul/mult_37_G2/ab[1][0] , \mat_mul/mult_37_G2/ab[1][1] ,
         \mat_mul/mult_37_G2/ab[1][2] , \mat_mul/mult_37_G2/ab[1][3] ,
         \mat_mul/mult_37_G2/ab[1][4] , \mat_mul/mult_37_G2/ab[1][5] ,
         \mat_mul/mult_37_G2/ab[1][6] , \mat_mul/mult_37_G2/ab[2][0] ,
         \mat_mul/mult_37_G2/ab[2][1] , \mat_mul/mult_37_G2/ab[2][2] ,
         \mat_mul/mult_37_G2/ab[2][3] , \mat_mul/mult_37_G2/ab[2][4] ,
         \mat_mul/mult_37_G2/ab[2][5] , \mat_mul/mult_37_G2/ab[3][0] ,
         \mat_mul/mult_37_G2/ab[3][1] , \mat_mul/mult_37_G2/ab[3][2] ,
         \mat_mul/mult_37_G2/ab[3][3] , \mat_mul/mult_37_G2/ab[3][4] ,
         \mat_mul/mult_37_G2/ab[4][0] , \mat_mul/mult_37_G2/ab[4][1] ,
         \mat_mul/mult_37_G2/ab[4][2] , \mat_mul/mult_37_G2/ab[4][3] ,
         \mat_mul/mult_37_G2/ab[5][0] , \mat_mul/mult_37_G2/ab[5][1] ,
         \mat_mul/mult_37_G2/ab[5][2] , \mat_mul/mult_37_G2/ab[6][0] ,
         \mat_mul/mult_37_G2/ab[6][1] , \mat_mul/mult_37_G2/ab[7][0] ,
         \mat_mul/mult_37_G2_G1_G2/FS_1/P[0][0][1] ,
         \mat_mul/mult_37_G2_G1_G2/FS_1/P[0][0][2] ,
         \mat_mul/mult_37_G2_G1_G2/FS_1/P[0][0][3] ,
         \mat_mul/mult_37_G2_G1_G2/FS_1/P[0][1][1] ,
         \mat_mul/mult_37_G2_G1_G2/FS_1/TEMP_P[0][0][0] ,
         \mat_mul/mult_37_G2_G1_G2/FS_1/TEMP_P[0][1][0] ,
         \mat_mul/mult_37_G2_G1_G2/A1[0] , \mat_mul/mult_37_G2_G1_G2/A1[1] ,
         \mat_mul/mult_37_G2_G1_G2/A1[2] , \mat_mul/mult_37_G2_G1_G2/A1[3] ,
         \mat_mul/mult_37_G2_G1_G2/A1[4] , \mat_mul/mult_37_G2_G1_G2/A1[5] ,
         \mat_mul/mult_37_G2_G1_G2/A_notx[0] ,
         \mat_mul/mult_37_G2_G1_G2/B_notx[0] ,
         \mat_mul/mult_37_G2_G1_G2/ab[0][1] ,
         \mat_mul/mult_37_G2_G1_G2/ab[0][2] ,
         \mat_mul/mult_37_G2_G1_G2/ab[0][3] ,
         \mat_mul/mult_37_G2_G1_G2/ab[0][4] ,
         \mat_mul/mult_37_G2_G1_G2/ab[0][5] ,
         \mat_mul/mult_37_G2_G1_G2/ab[0][6] ,
         \mat_mul/mult_37_G2_G1_G2/ab[0][7] ,
         \mat_mul/mult_37_G2_G1_G2/ab[1][0] ,
         \mat_mul/mult_37_G2_G1_G2/ab[1][1] ,
         \mat_mul/mult_37_G2_G1_G2/ab[1][2] ,
         \mat_mul/mult_37_G2_G1_G2/ab[1][3] ,
         \mat_mul/mult_37_G2_G1_G2/ab[1][4] ,
         \mat_mul/mult_37_G2_G1_G2/ab[1][5] ,
         \mat_mul/mult_37_G2_G1_G2/ab[1][6] ,
         \mat_mul/mult_37_G2_G1_G2/ab[2][0] ,
         \mat_mul/mult_37_G2_G1_G2/ab[2][1] ,
         \mat_mul/mult_37_G2_G1_G2/ab[2][2] ,
         \mat_mul/mult_37_G2_G1_G2/ab[2][3] ,
         \mat_mul/mult_37_G2_G1_G2/ab[2][4] ,
         \mat_mul/mult_37_G2_G1_G2/ab[2][5] ,
         \mat_mul/mult_37_G2_G1_G2/ab[3][0] ,
         \mat_mul/mult_37_G2_G1_G2/ab[3][1] ,
         \mat_mul/mult_37_G2_G1_G2/ab[3][2] ,
         \mat_mul/mult_37_G2_G1_G2/ab[3][3] ,
         \mat_mul/mult_37_G2_G1_G2/ab[3][4] ,
         \mat_mul/mult_37_G2_G1_G2/ab[4][0] ,
         \mat_mul/mult_37_G2_G1_G2/ab[4][1] ,
         \mat_mul/mult_37_G2_G1_G2/ab[4][2] ,
         \mat_mul/mult_37_G2_G1_G2/ab[4][3] ,
         \mat_mul/mult_37_G2_G1_G2/ab[5][0] ,
         \mat_mul/mult_37_G2_G1_G2/ab[5][1] ,
         \mat_mul/mult_37_G2_G1_G2/ab[5][2] ,
         \mat_mul/mult_37_G2_G1_G2/ab[6][0] ,
         \mat_mul/mult_37_G2_G1_G2/ab[6][1] ,
         \mat_mul/mult_37_G2_G1_G2/ab[7][0] ,
         \mat_mul/mult_37_G2_G2/FS_1/P[0][0][1] ,
         \mat_mul/mult_37_G2_G2/FS_1/P[0][0][2] ,
         \mat_mul/mult_37_G2_G2/FS_1/P[0][0][3] ,
         \mat_mul/mult_37_G2_G2/FS_1/P[0][1][1] ,
         \mat_mul/mult_37_G2_G2/FS_1/TEMP_P[0][0][0] ,
         \mat_mul/mult_37_G2_G2/FS_1/TEMP_P[0][1][0] ,
         \mat_mul/mult_37_G2_G2/A1[0] , \mat_mul/mult_37_G2_G2/A1[1] ,
         \mat_mul/mult_37_G2_G2/A1[2] , \mat_mul/mult_37_G2_G2/A1[3] ,
         \mat_mul/mult_37_G2_G2/A1[4] , \mat_mul/mult_37_G2_G2/A1[5] ,
         \mat_mul/mult_37_G2_G2/A_notx[0] , \mat_mul/mult_37_G2_G2/B_notx[0] ,
         \mat_mul/mult_37_G2_G2/ab[0][1] , \mat_mul/mult_37_G2_G2/ab[0][2] ,
         \mat_mul/mult_37_G2_G2/ab[0][3] , \mat_mul/mult_37_G2_G2/ab[0][4] ,
         \mat_mul/mult_37_G2_G2/ab[0][5] , \mat_mul/mult_37_G2_G2/ab[0][6] ,
         \mat_mul/mult_37_G2_G2/ab[0][7] , \mat_mul/mult_37_G2_G2/ab[1][0] ,
         \mat_mul/mult_37_G2_G2/ab[1][1] , \mat_mul/mult_37_G2_G2/ab[1][2] ,
         \mat_mul/mult_37_G2_G2/ab[1][3] , \mat_mul/mult_37_G2_G2/ab[1][4] ,
         \mat_mul/mult_37_G2_G2/ab[1][5] , \mat_mul/mult_37_G2_G2/ab[1][6] ,
         \mat_mul/mult_37_G2_G2/ab[2][0] , \mat_mul/mult_37_G2_G2/ab[2][1] ,
         \mat_mul/mult_37_G2_G2/ab[2][2] , \mat_mul/mult_37_G2_G2/ab[2][3] ,
         \mat_mul/mult_37_G2_G2/ab[2][4] , \mat_mul/mult_37_G2_G2/ab[2][5] ,
         \mat_mul/mult_37_G2_G2/ab[3][0] , \mat_mul/mult_37_G2_G2/ab[3][1] ,
         \mat_mul/mult_37_G2_G2/ab[3][2] , \mat_mul/mult_37_G2_G2/ab[3][3] ,
         \mat_mul/mult_37_G2_G2/ab[3][4] , \mat_mul/mult_37_G2_G2/ab[4][0] ,
         \mat_mul/mult_37_G2_G2/ab[4][1] , \mat_mul/mult_37_G2_G2/ab[4][2] ,
         \mat_mul/mult_37_G2_G2/ab[4][3] , \mat_mul/mult_37_G2_G2/ab[5][0] ,
         \mat_mul/mult_37_G2_G2/ab[5][1] , \mat_mul/mult_37_G2_G2/ab[5][2] ,
         \mat_mul/mult_37_G2_G2/ab[6][0] , \mat_mul/mult_37_G2_G2/ab[6][1] ,
         \mat_mul/mult_37_G2_G2/ab[7][0] ,
         \mat_mul/mult_37_G2_G2_G2/FS_1/P[0][0][1] ,
         \mat_mul/mult_37_G2_G2_G2/FS_1/P[0][0][2] ,
         \mat_mul/mult_37_G2_G2_G2/FS_1/P[0][0][3] ,
         \mat_mul/mult_37_G2_G2_G2/FS_1/P[0][1][1] ,
         \mat_mul/mult_37_G2_G2_G2/FS_1/TEMP_P[0][0][0] ,
         \mat_mul/mult_37_G2_G2_G2/FS_1/TEMP_P[0][1][0] ,
         \mat_mul/mult_37_G2_G2_G2/A1[0] , \mat_mul/mult_37_G2_G2_G2/A1[1] ,
         \mat_mul/mult_37_G2_G2_G2/A1[2] , \mat_mul/mult_37_G2_G2_G2/A1[3] ,
         \mat_mul/mult_37_G2_G2_G2/A1[4] , \mat_mul/mult_37_G2_G2_G2/A1[5] ,
         \mat_mul/mult_37_G2_G2_G2/A_notx[0] ,
         \mat_mul/mult_37_G2_G2_G2/B_notx[0] ,
         \mat_mul/mult_37_G2_G2_G2/ab[0][1] ,
         \mat_mul/mult_37_G2_G2_G2/ab[0][2] ,
         \mat_mul/mult_37_G2_G2_G2/ab[0][3] ,
         \mat_mul/mult_37_G2_G2_G2/ab[0][4] ,
         \mat_mul/mult_37_G2_G2_G2/ab[0][5] ,
         \mat_mul/mult_37_G2_G2_G2/ab[0][6] ,
         \mat_mul/mult_37_G2_G2_G2/ab[0][7] ,
         \mat_mul/mult_37_G2_G2_G2/ab[1][0] ,
         \mat_mul/mult_37_G2_G2_G2/ab[1][1] ,
         \mat_mul/mult_37_G2_G2_G2/ab[1][2] ,
         \mat_mul/mult_37_G2_G2_G2/ab[1][3] ,
         \mat_mul/mult_37_G2_G2_G2/ab[1][4] ,
         \mat_mul/mult_37_G2_G2_G2/ab[1][5] ,
         \mat_mul/mult_37_G2_G2_G2/ab[1][6] ,
         \mat_mul/mult_37_G2_G2_G2/ab[2][0] ,
         \mat_mul/mult_37_G2_G2_G2/ab[2][1] ,
         \mat_mul/mult_37_G2_G2_G2/ab[2][2] ,
         \mat_mul/mult_37_G2_G2_G2/ab[2][3] ,
         \mat_mul/mult_37_G2_G2_G2/ab[2][4] ,
         \mat_mul/mult_37_G2_G2_G2/ab[2][5] ,
         \mat_mul/mult_37_G2_G2_G2/ab[3][0] ,
         \mat_mul/mult_37_G2_G2_G2/ab[3][1] ,
         \mat_mul/mult_37_G2_G2_G2/ab[3][2] ,
         \mat_mul/mult_37_G2_G2_G2/ab[3][3] ,
         \mat_mul/mult_37_G2_G2_G2/ab[3][4] ,
         \mat_mul/mult_37_G2_G2_G2/ab[4][0] ,
         \mat_mul/mult_37_G2_G2_G2/ab[4][1] ,
         \mat_mul/mult_37_G2_G2_G2/ab[4][2] ,
         \mat_mul/mult_37_G2_G2_G2/ab[4][3] ,
         \mat_mul/mult_37_G2_G2_G2/ab[5][0] ,
         \mat_mul/mult_37_G2_G2_G2/ab[5][1] ,
         \mat_mul/mult_37_G2_G2_G2/ab[5][2] ,
         \mat_mul/mult_37_G2_G2_G2/ab[6][0] ,
         \mat_mul/mult_37_G2_G2_G2/ab[6][1] ,
         \mat_mul/mult_37_G2_G2_G2/ab[7][0] , n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413;
  wire   [31:0] m_add;
  wire   [31:0] m_sub;
  wire   [31:0] m_mul;
  wire   [127:0] m_kro;
  wire   [7:0] \mat_sub/r106/B_AS ;
  wire   [7:0] \mat_sub/r94/B_AS ;
  wire   [7:0] \mat_sub/r102/B_AS ;
  wire   [7:0] \mat_sub/r98/B_AS ;
  wire   [7:0] \mat_kron/mult_40/B_not ;
  wire   [7:0] \mat_kron/mult_40/A_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G1_G1_G1/B_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G1_G1_G1/A_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G1_G1/B_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G1_G1/A_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G2_G1_G1/B_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G2_G1_G1/A_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G1/B_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G1/A_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G1_G2_G1/B_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G1_G2_G1/A_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G2_G1/B_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G2_G1/A_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G2_G2_G1/B_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G2_G2_G1/A_not ;
  wire   [7:0] \mat_kron/mult_40_G2/B_not ;
  wire   [7:0] \mat_kron/mult_40_G2/A_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G1_G1_G2/B_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G1_G1_G2/A_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G1_G2/B_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G1_G2/A_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G2_G1_G2/B_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G2_G1_G2/A_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G2/B_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G2/A_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G1_G2_G2/B_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G1_G2_G2/A_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G2_G2/B_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G2_G2/A_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G2_G2_G2/B_not ;
  wire   [7:0] \mat_kron/mult_40_G2_G2_G2_G2/A_not ;
  wire   [7:0] \mat_mul/mult_37/B_not ;
  wire   [7:0] \mat_mul/mult_37/A_not ;
  wire   [7:0] \mat_mul/mult_37_G2_G1_G1/B_not ;
  wire   [7:0] \mat_mul/mult_37_G2_G1_G1/A_not ;
  wire   [7:0] \mat_mul/mult_37_G2_G1/B_not ;
  wire   [7:0] \mat_mul/mult_37_G2_G1/A_not ;
  wire   [7:0] \mat_mul/mult_37_G2_G2_G1/B_not ;
  wire   [7:0] \mat_mul/mult_37_G2_G2_G1/A_not ;
  wire   [7:0] \mat_mul/mult_37_G2/B_not ;
  wire   [7:0] \mat_mul/mult_37_G2/A_not ;
  wire   [7:0] \mat_mul/mult_37_G2_G1_G2/B_not ;
  wire   [7:0] \mat_mul/mult_37_G2_G1_G2/A_not ;
  wire   [7:0] \mat_mul/mult_37_G2_G2/B_not ;
  wire   [7:0] \mat_mul/mult_37_G2_G2/A_not ;
  wire   [7:0] \mat_mul/mult_37_G2_G2_G2/B_not ;
  wire   [7:0] \mat_mul/mult_37_G2_G2_G2/A_not ;
  wire   [7:0] \mat_add/r106/B_AS ;
  wire   [7:0] \mat_add/r94/B_AS ;
  wire   [7:0] \mat_add/r102/B_AS ;
  wire   [7:0] \mat_add/r98/B_AS ;
  assign \mat_add/r106/B_AS  [7] = B[7];
  assign \mat_add/r106/B_AS  [6] = B[6];
  assign \mat_add/r106/B_AS  [5] = B[5];
  assign \mat_add/r106/B_AS  [4] = B[4];
  assign \mat_add/r106/B_AS  [3] = B[3];
  assign \mat_add/r106/B_AS  [2] = B[2];
  assign \mat_add/r106/B_AS  [1] = B[1];
  assign \mat_add/r106/B_AS  [0] = B[0];
  assign \mat_add/r94/B_AS  [7] = B[31];
  assign \mat_add/r94/B_AS  [6] = B[30];
  assign \mat_add/r94/B_AS  [5] = B[29];
  assign \mat_add/r94/B_AS  [4] = B[28];
  assign \mat_add/r94/B_AS  [3] = B[27];
  assign \mat_add/r94/B_AS  [2] = B[26];
  assign \mat_add/r94/B_AS  [1] = B[25];
  assign \mat_add/r94/B_AS  [0] = B[24];
  assign \mat_add/r102/B_AS  [7] = B[15];
  assign \mat_add/r102/B_AS  [6] = B[14];
  assign \mat_add/r102/B_AS  [5] = B[13];
  assign \mat_add/r102/B_AS  [4] = B[12];
  assign \mat_add/r102/B_AS  [3] = B[11];
  assign \mat_add/r102/B_AS  [2] = B[10];
  assign \mat_add/r102/B_AS  [1] = B[9];
  assign \mat_add/r102/B_AS  [0] = B[8];
  assign \mat_add/r98/B_AS  [7] = B[23];
  assign \mat_add/r98/B_AS  [6] = B[22];
  assign \mat_add/r98/B_AS  [5] = B[21];
  assign \mat_add/r98/B_AS  [4] = B[20];
  assign \mat_add/r98/B_AS  [3] = B[19];
  assign \mat_add/r98/B_AS  [2] = B[18];
  assign \mat_add/r98/B_AS  [1] = B[17];
  assign \mat_add/r98/B_AS  [0] = B[16];

  nand2 C410 ( .a(op[0]), .b(op[1]), .out(n1) );
  inv I_4 ( .in(N139), .out(N140) );
  nand2 C408 ( .a(N135), .b(op[1]), .out(N139) );
  inv I_2 ( .in(N136), .out(N137) );
  nand2 C405 ( .a(op[0]), .b(n163), .out(N136) );
  inv I_1 ( .in(op[0]), .out(N135) );
  inv I_0 ( .in(N133), .out(N134) );
  nand2 C402 ( .a(N135), .b(n163), .out(N133) );
  dff \C_reg_reg[127]  ( .d(N132), .gclk(clk), .rnot(resetn), .q(C[127]) );
  dff \C_reg_reg[126]  ( .d(N131), .gclk(clk), .rnot(resetn), .q(C[126]) );
  dff \C_reg_reg[125]  ( .d(N130), .gclk(clk), .rnot(resetn), .q(C[125]) );
  dff \C_reg_reg[124]  ( .d(N129), .gclk(clk), .rnot(resetn), .q(C[124]) );
  dff \C_reg_reg[123]  ( .d(N128), .gclk(clk), .rnot(resetn), .q(C[123]) );
  dff \C_reg_reg[122]  ( .d(N127), .gclk(clk), .rnot(resetn), .q(C[122]) );
  dff \C_reg_reg[121]  ( .d(N126), .gclk(clk), .rnot(resetn), .q(C[121]) );
  dff \C_reg_reg[120]  ( .d(N125), .gclk(clk), .rnot(resetn), .q(C[120]) );
  dff \C_reg_reg[119]  ( .d(N124), .gclk(clk), .rnot(resetn), .q(C[119]) );
  dff \C_reg_reg[118]  ( .d(N123), .gclk(clk), .rnot(resetn), .q(C[118]) );
  dff \C_reg_reg[117]  ( .d(N122), .gclk(clk), .rnot(resetn), .q(C[117]) );
  dff \C_reg_reg[116]  ( .d(N121), .gclk(clk), .rnot(resetn), .q(C[116]) );
  dff \C_reg_reg[115]  ( .d(N120), .gclk(clk), .rnot(resetn), .q(C[115]) );
  dff \C_reg_reg[114]  ( .d(N119), .gclk(clk), .rnot(resetn), .q(C[114]) );
  dff \C_reg_reg[113]  ( .d(N118), .gclk(clk), .rnot(resetn), .q(C[113]) );
  dff \C_reg_reg[112]  ( .d(N117), .gclk(clk), .rnot(resetn), .q(C[112]) );
  dff \C_reg_reg[111]  ( .d(N116), .gclk(clk), .rnot(resetn), .q(C[111]) );
  dff \C_reg_reg[110]  ( .d(N115), .gclk(clk), .rnot(resetn), .q(C[110]) );
  dff \C_reg_reg[109]  ( .d(N114), .gclk(clk), .rnot(resetn), .q(C[109]) );
  dff \C_reg_reg[108]  ( .d(N113), .gclk(clk), .rnot(resetn), .q(C[108]) );
  dff \C_reg_reg[107]  ( .d(N112), .gclk(clk), .rnot(resetn), .q(C[107]) );
  dff \C_reg_reg[106]  ( .d(N111), .gclk(clk), .rnot(resetn), .q(C[106]) );
  dff \C_reg_reg[105]  ( .d(N110), .gclk(clk), .rnot(resetn), .q(C[105]) );
  dff \C_reg_reg[104]  ( .d(N109), .gclk(clk), .rnot(resetn), .q(C[104]) );
  dff \C_reg_reg[103]  ( .d(N108), .gclk(clk), .rnot(resetn), .q(C[103]) );
  dff \C_reg_reg[102]  ( .d(N107), .gclk(clk), .rnot(resetn), .q(C[102]) );
  dff \C_reg_reg[101]  ( .d(N106), .gclk(clk), .rnot(resetn), .q(C[101]) );
  dff \C_reg_reg[100]  ( .d(N105), .gclk(clk), .rnot(resetn), .q(C[100]) );
  dff \C_reg_reg[99]  ( .d(N104), .gclk(clk), .rnot(resetn), .q(C[99]) );
  dff \C_reg_reg[98]  ( .d(N103), .gclk(clk), .rnot(resetn), .q(C[98]) );
  dff \C_reg_reg[97]  ( .d(N102), .gclk(clk), .rnot(resetn), .q(C[97]) );
  dff \C_reg_reg[96]  ( .d(N101), .gclk(clk), .rnot(resetn), .q(C[96]) );
  dff \C_reg_reg[95]  ( .d(N100), .gclk(clk), .rnot(resetn), .q(C[95]) );
  dff \C_reg_reg[94]  ( .d(N99), .gclk(clk), .rnot(resetn), .q(C[94]) );
  dff \C_reg_reg[93]  ( .d(N98), .gclk(clk), .rnot(resetn), .q(C[93]) );
  dff \C_reg_reg[92]  ( .d(N97), .gclk(clk), .rnot(resetn), .q(C[92]) );
  dff \C_reg_reg[91]  ( .d(N96), .gclk(clk), .rnot(resetn), .q(C[91]) );
  dff \C_reg_reg[90]  ( .d(N95), .gclk(clk), .rnot(resetn), .q(C[90]) );
  dff \C_reg_reg[89]  ( .d(N94), .gclk(clk), .rnot(resetn), .q(C[89]) );
  dff \C_reg_reg[88]  ( .d(N93), .gclk(clk), .rnot(resetn), .q(C[88]) );
  dff \C_reg_reg[87]  ( .d(N92), .gclk(clk), .rnot(resetn), .q(C[87]) );
  dff \C_reg_reg[86]  ( .d(N91), .gclk(clk), .rnot(resetn), .q(C[86]) );
  dff \C_reg_reg[85]  ( .d(N90), .gclk(clk), .rnot(resetn), .q(C[85]) );
  dff \C_reg_reg[84]  ( .d(N89), .gclk(clk), .rnot(resetn), .q(C[84]) );
  dff \C_reg_reg[83]  ( .d(N88), .gclk(clk), .rnot(resetn), .q(C[83]) );
  dff \C_reg_reg[82]  ( .d(N87), .gclk(clk), .rnot(resetn), .q(C[82]) );
  dff \C_reg_reg[81]  ( .d(N86), .gclk(clk), .rnot(resetn), .q(C[81]) );
  dff \C_reg_reg[80]  ( .d(N85), .gclk(clk), .rnot(resetn), .q(C[80]) );
  dff \C_reg_reg[79]  ( .d(N84), .gclk(clk), .rnot(resetn), .q(C[79]) );
  dff \C_reg_reg[78]  ( .d(N83), .gclk(clk), .rnot(resetn), .q(C[78]) );
  dff \C_reg_reg[77]  ( .d(N82), .gclk(clk), .rnot(resetn), .q(C[77]) );
  dff \C_reg_reg[76]  ( .d(N81), .gclk(clk), .rnot(resetn), .q(C[76]) );
  dff \C_reg_reg[75]  ( .d(N80), .gclk(clk), .rnot(resetn), .q(C[75]) );
  dff \C_reg_reg[74]  ( .d(N79), .gclk(clk), .rnot(resetn), .q(C[74]) );
  dff \C_reg_reg[73]  ( .d(N78), .gclk(clk), .rnot(resetn), .q(C[73]) );
  dff \C_reg_reg[72]  ( .d(N77), .gclk(clk), .rnot(resetn), .q(C[72]) );
  dff \C_reg_reg[71]  ( .d(N76), .gclk(clk), .rnot(resetn), .q(C[71]) );
  dff \C_reg_reg[70]  ( .d(N75), .gclk(clk), .rnot(resetn), .q(C[70]) );
  dff \C_reg_reg[69]  ( .d(N74), .gclk(clk), .rnot(resetn), .q(C[69]) );
  dff \C_reg_reg[68]  ( .d(N73), .gclk(clk), .rnot(resetn), .q(C[68]) );
  dff \C_reg_reg[67]  ( .d(N72), .gclk(clk), .rnot(resetn), .q(C[67]) );
  dff \C_reg_reg[66]  ( .d(N71), .gclk(clk), .rnot(resetn), .q(C[66]) );
  dff \C_reg_reg[65]  ( .d(N70), .gclk(clk), .rnot(resetn), .q(C[65]) );
  dff \C_reg_reg[64]  ( .d(N69), .gclk(clk), .rnot(resetn), .q(C[64]) );
  dff \C_reg_reg[63]  ( .d(N68), .gclk(clk), .rnot(resetn), .q(C[63]) );
  dff \C_reg_reg[62]  ( .d(N67), .gclk(clk), .rnot(resetn), .q(C[62]) );
  dff \C_reg_reg[61]  ( .d(N66), .gclk(clk), .rnot(resetn), .q(C[61]) );
  dff \C_reg_reg[60]  ( .d(N65), .gclk(clk), .rnot(resetn), .q(C[60]) );
  dff \C_reg_reg[59]  ( .d(N64), .gclk(clk), .rnot(resetn), .q(C[59]) );
  dff \C_reg_reg[58]  ( .d(N63), .gclk(clk), .rnot(resetn), .q(C[58]) );
  dff \C_reg_reg[57]  ( .d(N62), .gclk(clk), .rnot(resetn), .q(C[57]) );
  dff \C_reg_reg[56]  ( .d(N61), .gclk(clk), .rnot(resetn), .q(C[56]) );
  dff \C_reg_reg[55]  ( .d(N60), .gclk(clk), .rnot(resetn), .q(C[55]) );
  dff \C_reg_reg[54]  ( .d(N59), .gclk(clk), .rnot(resetn), .q(C[54]) );
  dff \C_reg_reg[53]  ( .d(N58), .gclk(clk), .rnot(resetn), .q(C[53]) );
  dff \C_reg_reg[52]  ( .d(N57), .gclk(clk), .rnot(resetn), .q(C[52]) );
  dff \C_reg_reg[51]  ( .d(N56), .gclk(clk), .rnot(resetn), .q(C[51]) );
  dff \C_reg_reg[50]  ( .d(N55), .gclk(clk), .rnot(resetn), .q(C[50]) );
  dff \C_reg_reg[49]  ( .d(N54), .gclk(clk), .rnot(resetn), .q(C[49]) );
  dff \C_reg_reg[48]  ( .d(N53), .gclk(clk), .rnot(resetn), .q(C[48]) );
  dff \C_reg_reg[47]  ( .d(N52), .gclk(clk), .rnot(resetn), .q(C[47]) );
  dff \C_reg_reg[46]  ( .d(N51), .gclk(clk), .rnot(resetn), .q(C[46]) );
  dff \C_reg_reg[45]  ( .d(N50), .gclk(clk), .rnot(resetn), .q(C[45]) );
  dff \C_reg_reg[44]  ( .d(N49), .gclk(clk), .rnot(resetn), .q(C[44]) );
  dff \C_reg_reg[43]  ( .d(N48), .gclk(clk), .rnot(resetn), .q(C[43]) );
  dff \C_reg_reg[42]  ( .d(N47), .gclk(clk), .rnot(resetn), .q(C[42]) );
  dff \C_reg_reg[41]  ( .d(N46), .gclk(clk), .rnot(resetn), .q(C[41]) );
  dff \C_reg_reg[40]  ( .d(N45), .gclk(clk), .rnot(resetn), .q(C[40]) );
  dff \C_reg_reg[39]  ( .d(N44), .gclk(clk), .rnot(resetn), .q(C[39]) );
  dff \C_reg_reg[38]  ( .d(N43), .gclk(clk), .rnot(resetn), .q(C[38]) );
  dff \C_reg_reg[37]  ( .d(N42), .gclk(clk), .rnot(resetn), .q(C[37]) );
  dff \C_reg_reg[36]  ( .d(N41), .gclk(clk), .rnot(resetn), .q(C[36]) );
  dff \C_reg_reg[35]  ( .d(N40), .gclk(clk), .rnot(resetn), .q(C[35]) );
  dff \C_reg_reg[34]  ( .d(N39), .gclk(clk), .rnot(resetn), .q(C[34]) );
  dff \C_reg_reg[33]  ( .d(N38), .gclk(clk), .rnot(resetn), .q(C[33]) );
  dff \C_reg_reg[32]  ( .d(N37), .gclk(clk), .rnot(resetn), .q(C[32]) );
  dff \C_reg_reg[31]  ( .d(N36), .gclk(clk), .rnot(resetn), .q(C[31]) );
  dff \C_reg_reg[30]  ( .d(N35), .gclk(clk), .rnot(resetn), .q(C[30]) );
  dff \C_reg_reg[29]  ( .d(N34), .gclk(clk), .rnot(resetn), .q(C[29]) );
  dff \C_reg_reg[28]  ( .d(N33), .gclk(clk), .rnot(resetn), .q(C[28]) );
  dff \C_reg_reg[27]  ( .d(N32), .gclk(clk), .rnot(resetn), .q(C[27]) );
  dff \C_reg_reg[26]  ( .d(N31), .gclk(clk), .rnot(resetn), .q(C[26]) );
  dff \C_reg_reg[25]  ( .d(N30), .gclk(clk), .rnot(resetn), .q(C[25]) );
  dff \C_reg_reg[24]  ( .d(N29), .gclk(clk), .rnot(resetn), .q(C[24]) );
  dff \C_reg_reg[23]  ( .d(N28), .gclk(clk), .rnot(resetn), .q(C[23]) );
  dff \C_reg_reg[22]  ( .d(N27), .gclk(clk), .rnot(resetn), .q(C[22]) );
  dff \C_reg_reg[21]  ( .d(N26), .gclk(clk), .rnot(resetn), .q(C[21]) );
  dff \C_reg_reg[20]  ( .d(N25), .gclk(clk), .rnot(resetn), .q(C[20]) );
  dff \C_reg_reg[19]  ( .d(N24), .gclk(clk), .rnot(resetn), .q(C[19]) );
  dff \C_reg_reg[18]  ( .d(N23), .gclk(clk), .rnot(resetn), .q(C[18]) );
  dff \C_reg_reg[17]  ( .d(N22), .gclk(clk), .rnot(resetn), .q(C[17]) );
  dff \C_reg_reg[16]  ( .d(N21), .gclk(clk), .rnot(resetn), .q(C[16]) );
  dff \C_reg_reg[15]  ( .d(N20), .gclk(clk), .rnot(resetn), .q(C[15]) );
  dff \C_reg_reg[14]  ( .d(N19), .gclk(clk), .rnot(resetn), .q(C[14]) );
  dff \C_reg_reg[13]  ( .d(N18), .gclk(clk), .rnot(resetn), .q(C[13]) );
  dff \C_reg_reg[12]  ( .d(N17), .gclk(clk), .rnot(resetn), .q(C[12]) );
  dff \C_reg_reg[11]  ( .d(N16), .gclk(clk), .rnot(resetn), .q(C[11]) );
  dff \C_reg_reg[10]  ( .d(N15), .gclk(clk), .rnot(resetn), .q(C[10]) );
  dff \C_reg_reg[9]  ( .d(N14), .gclk(clk), .rnot(resetn), .q(C[9]) );
  dff \C_reg_reg[8]  ( .d(N13), .gclk(clk), .rnot(resetn), .q(C[8]) );
  dff \C_reg_reg[7]  ( .d(N12), .gclk(clk), .rnot(resetn), .q(C[7]) );
  dff \C_reg_reg[6]  ( .d(N11), .gclk(clk), .rnot(resetn), .q(C[6]) );
  dff \C_reg_reg[5]  ( .d(N10), .gclk(clk), .rnot(resetn), .q(C[5]) );
  dff \C_reg_reg[4]  ( .d(N9), .gclk(clk), .rnot(resetn), .q(C[4]) );
  dff \C_reg_reg[3]  ( .d(N8), .gclk(clk), .rnot(resetn), .q(C[3]) );
  dff \C_reg_reg[2]  ( .d(N7), .gclk(clk), .rnot(resetn), .q(C[2]) );
  dff \C_reg_reg[1]  ( .d(N6), .gclk(clk), .rnot(resetn), .q(C[1]) );
  dff \C_reg_reg[0]  ( .d(N5), .gclk(clk), .rnot(resetn), .q(C[0]) );
  nor2 U3 ( .a(n1), .b(n2), .out(N99) );
  inv U4 ( .in(m_kro[94]), .out(n2) );
  nor2 U5 ( .a(n1), .b(n3), .out(N98) );
  inv U6 ( .in(m_kro[93]), .out(n3) );
  nor2 U7 ( .a(n1), .b(n4), .out(N97) );
  inv U8 ( .in(m_kro[92]), .out(n4) );
  nor2 U9 ( .a(n1), .b(n5), .out(N96) );
  inv U10 ( .in(m_kro[91]), .out(n5) );
  nor2 U11 ( .a(n1), .b(n6), .out(N95) );
  inv U12 ( .in(m_kro[90]), .out(n6) );
  nor2 U13 ( .a(n1), .b(n7), .out(N94) );
  inv U14 ( .in(m_kro[89]), .out(n7) );
  nor2 U15 ( .a(n1), .b(n8), .out(N93) );
  inv U16 ( .in(m_kro[88]), .out(n8) );
  nor2 U17 ( .a(n1), .b(n9), .out(N92) );
  inv U18 ( .in(m_kro[87]), .out(n9) );
  nor2 U19 ( .a(n1), .b(n10), .out(N91) );
  inv U20 ( .in(m_kro[86]), .out(n10) );
  nor2 U21 ( .a(n1), .b(n11), .out(N90) );
  inv U22 ( .in(m_kro[85]), .out(n11) );
  nand2 U23 ( .a(n12), .b(n13), .out(N9) );
  aoi22 U24 ( .a(m_add[4]), .b(N134), .c(m_sub[4]), .d(N137), .out(n13) );
  aoi22 U25 ( .a(m_mul[4]), .b(N140), .c(m_kro[4]), .d(n14), .out(n12) );
  nor2 U26 ( .a(n1), .b(n15), .out(N89) );
  inv U27 ( .in(m_kro[84]), .out(n15) );
  nor2 U28 ( .a(n1), .b(n16), .out(N88) );
  inv U29 ( .in(m_kro[83]), .out(n16) );
  nor2 U30 ( .a(n1), .b(n17), .out(N87) );
  inv U31 ( .in(m_kro[82]), .out(n17) );
  nor2 U32 ( .a(n1), .b(n18), .out(N86) );
  inv U33 ( .in(m_kro[81]), .out(n18) );
  nor2 U34 ( .a(n1), .b(n19), .out(N85) );
  inv U35 ( .in(m_kro[80]), .out(n19) );
  nor2 U36 ( .a(n1), .b(n20), .out(N84) );
  inv U37 ( .in(m_kro[79]), .out(n20) );
  nor2 U38 ( .a(n1), .b(n21), .out(N83) );
  inv U39 ( .in(m_kro[78]), .out(n21) );
  nor2 U40 ( .a(n1), .b(n22), .out(N82) );
  inv U41 ( .in(m_kro[77]), .out(n22) );
  nor2 U42 ( .a(n1), .b(n23), .out(N81) );
  inv U43 ( .in(m_kro[76]), .out(n23) );
  nor2 U44 ( .a(n1), .b(n24), .out(N80) );
  inv U45 ( .in(m_kro[75]), .out(n24) );
  nand2 U46 ( .a(n25), .b(n26), .out(N8) );
  aoi22 U47 ( .a(m_add[3]), .b(N134), .c(m_sub[3]), .d(N137), .out(n26) );
  aoi22 U48 ( .a(m_mul[3]), .b(N140), .c(m_kro[3]), .d(n14), .out(n25) );
  nor2 U49 ( .a(n1), .b(n27), .out(N79) );
  inv U50 ( .in(m_kro[74]), .out(n27) );
  nor2 U51 ( .a(n1), .b(n28), .out(N78) );
  inv U52 ( .in(m_kro[73]), .out(n28) );
  nor2 U53 ( .a(n1), .b(n29), .out(N77) );
  inv U54 ( .in(m_kro[72]), .out(n29) );
  nor2 U55 ( .a(n1), .b(n30), .out(N76) );
  inv U56 ( .in(m_kro[71]), .out(n30) );
  nor2 U57 ( .a(n1), .b(n31), .out(N75) );
  inv U58 ( .in(m_kro[70]), .out(n31) );
  nor2 U59 ( .a(n1), .b(n32), .out(N74) );
  inv U60 ( .in(m_kro[69]), .out(n32) );
  nor2 U61 ( .a(n1), .b(n33), .out(N73) );
  inv U62 ( .in(m_kro[68]), .out(n33) );
  nor2 U63 ( .a(n1), .b(n34), .out(N72) );
  inv U64 ( .in(m_kro[67]), .out(n34) );
  nor2 U65 ( .a(n1), .b(n35), .out(N71) );
  inv U66 ( .in(m_kro[66]), .out(n35) );
  nor2 U67 ( .a(n1), .b(n36), .out(N70) );
  inv U68 ( .in(m_kro[65]), .out(n36) );
  nand2 U69 ( .a(n37), .b(n38), .out(N7) );
  aoi22 U70 ( .a(m_add[2]), .b(N134), .c(m_sub[2]), .d(N137), .out(n38) );
  aoi22 U71 ( .a(m_mul[2]), .b(N140), .c(m_kro[2]), .d(n14), .out(n37) );
  nor2 U72 ( .a(n1), .b(n39), .out(N69) );
  inv U73 ( .in(m_kro[64]), .out(n39) );
  nor2 U74 ( .a(n1), .b(n40), .out(N68) );
  inv U75 ( .in(m_kro[63]), .out(n40) );
  nor2 U76 ( .a(n1), .b(n41), .out(N67) );
  inv U77 ( .in(m_kro[62]), .out(n41) );
  nor2 U78 ( .a(n1), .b(n42), .out(N66) );
  inv U79 ( .in(m_kro[61]), .out(n42) );
  nor2 U80 ( .a(n1), .b(n43), .out(N65) );
  inv U81 ( .in(m_kro[60]), .out(n43) );
  nor2 U82 ( .a(n1), .b(n44), .out(N64) );
  inv U83 ( .in(m_kro[59]), .out(n44) );
  nor2 U84 ( .a(n1), .b(n45), .out(N63) );
  inv U85 ( .in(m_kro[58]), .out(n45) );
  nor2 U86 ( .a(n1), .b(n46), .out(N62) );
  inv U87 ( .in(m_kro[57]), .out(n46) );
  nor2 U88 ( .a(n1), .b(n47), .out(N61) );
  inv U89 ( .in(m_kro[56]), .out(n47) );
  nor2 U90 ( .a(n1), .b(n48), .out(N60) );
  inv U91 ( .in(m_kro[55]), .out(n48) );
  nand2 U92 ( .a(n49), .b(n50), .out(N6) );
  aoi22 U93 ( .a(m_add[1]), .b(N134), .c(m_sub[1]), .d(N137), .out(n50) );
  aoi22 U94 ( .a(m_mul[1]), .b(N140), .c(m_kro[1]), .d(n14), .out(n49) );
  nor2 U95 ( .a(n1), .b(n51), .out(N59) );
  inv U96 ( .in(m_kro[54]), .out(n51) );
  nor2 U97 ( .a(n1), .b(n52), .out(N58) );
  inv U98 ( .in(m_kro[53]), .out(n52) );
  nor2 U99 ( .a(n1), .b(n53), .out(N57) );
  inv U100 ( .in(m_kro[52]), .out(n53) );
  nor2 U101 ( .a(n1), .b(n54), .out(N56) );
  inv U102 ( .in(m_kro[51]), .out(n54) );
  nor2 U103 ( .a(n1), .b(n55), .out(N55) );
  inv U104 ( .in(m_kro[50]), .out(n55) );
  nor2 U105 ( .a(n1), .b(n56), .out(N54) );
  inv U106 ( .in(m_kro[49]), .out(n56) );
  nor2 U107 ( .a(n1), .b(n57), .out(N53) );
  inv U108 ( .in(m_kro[48]), .out(n57) );
  nor2 U109 ( .a(n1), .b(n58), .out(N52) );
  inv U110 ( .in(m_kro[47]), .out(n58) );
  nor2 U111 ( .a(n1), .b(n59), .out(N51) );
  inv U112 ( .in(m_kro[46]), .out(n59) );
  nor2 U113 ( .a(n1), .b(n60), .out(N50) );
  inv U114 ( .in(m_kro[45]), .out(n60) );
  nand2 U115 ( .a(n61), .b(n62), .out(N5) );
  aoi22 U116 ( .a(m_add[0]), .b(N134), .c(m_sub[0]), .d(N137), .out(n62) );
  aoi22 U117 ( .a(m_mul[0]), .b(N140), .c(m_kro[0]), .d(n14), .out(n61) );
  nor2 U118 ( .a(n1), .b(n63), .out(N49) );
  inv U119 ( .in(m_kro[44]), .out(n63) );
  nor2 U120 ( .a(n1), .b(n64), .out(N48) );
  inv U121 ( .in(m_kro[43]), .out(n64) );
  nor2 U122 ( .a(n1), .b(n65), .out(N47) );
  inv U123 ( .in(m_kro[42]), .out(n65) );
  nor2 U124 ( .a(n1), .b(n66), .out(N46) );
  inv U125 ( .in(m_kro[41]), .out(n66) );
  nor2 U126 ( .a(n1), .b(n67), .out(N45) );
  inv U127 ( .in(m_kro[40]), .out(n67) );
  nor2 U128 ( .a(n1), .b(n68), .out(N44) );
  inv U129 ( .in(m_kro[39]), .out(n68) );
  nor2 U130 ( .a(n1), .b(n69), .out(N43) );
  inv U131 ( .in(m_kro[38]), .out(n69) );
  nor2 U132 ( .a(n1), .b(n70), .out(N42) );
  inv U133 ( .in(m_kro[37]), .out(n70) );
  nor2 U134 ( .a(n1), .b(n71), .out(N41) );
  inv U135 ( .in(m_kro[36]), .out(n71) );
  nor2 U136 ( .a(n1), .b(n72), .out(N40) );
  inv U137 ( .in(m_kro[35]), .out(n72) );
  nor2 U138 ( .a(n1), .b(n73), .out(N39) );
  inv U139 ( .in(m_kro[34]), .out(n73) );
  nor2 U140 ( .a(n1), .b(n74), .out(N38) );
  inv U141 ( .in(m_kro[33]), .out(n74) );
  nor2 U142 ( .a(n1), .b(n75), .out(N37) );
  inv U143 ( .in(m_kro[32]), .out(n75) );
  nand2 U144 ( .a(n76), .b(n77), .out(N36) );
  aoi22 U145 ( .a(m_add[31]), .b(N134), .c(m_sub[31]), .d(N137), .out(n77) );
  aoi22 U146 ( .a(m_mul[31]), .b(N140), .c(m_kro[31]), .d(n14), .out(n76) );
  nand2 U147 ( .a(n78), .b(n79), .out(N35) );
  aoi22 U148 ( .a(m_add[30]), .b(N134), .c(m_sub[30]), .d(N137), .out(n79) );
  aoi22 U149 ( .a(m_mul[30]), .b(N140), .c(m_kro[30]), .d(n14), .out(n78) );
  nand2 U150 ( .a(n80), .b(n81), .out(N34) );
  aoi22 U151 ( .a(m_add[29]), .b(N134), .c(m_sub[29]), .d(N137), .out(n81) );
  aoi22 U152 ( .a(m_mul[29]), .b(N140), .c(m_kro[29]), .d(n14), .out(n80) );
  nand2 U153 ( .a(n82), .b(n83), .out(N33) );
  aoi22 U154 ( .a(m_add[28]), .b(N134), .c(m_sub[28]), .d(N137), .out(n83) );
  aoi22 U155 ( .a(m_mul[28]), .b(N140), .c(m_kro[28]), .d(n14), .out(n82) );
  nand2 U156 ( .a(n84), .b(n85), .out(N32) );
  aoi22 U157 ( .a(m_add[27]), .b(N134), .c(m_sub[27]), .d(N137), .out(n85) );
  aoi22 U158 ( .a(m_mul[27]), .b(N140), .c(m_kro[27]), .d(n14), .out(n84) );
  nand2 U159 ( .a(n86), .b(n87), .out(N31) );
  aoi22 U160 ( .a(m_add[26]), .b(N134), .c(m_sub[26]), .d(N137), .out(n87) );
  aoi22 U161 ( .a(m_mul[26]), .b(N140), .c(m_kro[26]), .d(n14), .out(n86) );
  nand2 U162 ( .a(n88), .b(n89), .out(N30) );
  aoi22 U163 ( .a(m_add[25]), .b(N134), .c(m_sub[25]), .d(N137), .out(n89) );
  aoi22 U164 ( .a(m_mul[25]), .b(N140), .c(m_kro[25]), .d(n14), .out(n88) );
  nand2 U165 ( .a(n90), .b(n91), .out(N29) );
  aoi22 U166 ( .a(m_add[24]), .b(N134), .c(m_sub[24]), .d(N137), .out(n91) );
  aoi22 U167 ( .a(m_mul[24]), .b(N140), .c(m_kro[24]), .d(n14), .out(n90) );
  nand2 U168 ( .a(n92), .b(n93), .out(N28) );
  aoi22 U169 ( .a(m_add[23]), .b(N134), .c(m_sub[23]), .d(N137), .out(n93) );
  aoi22 U170 ( .a(m_mul[23]), .b(N140), .c(m_kro[23]), .d(n14), .out(n92) );
  nand2 U171 ( .a(n94), .b(n95), .out(N27) );
  aoi22 U172 ( .a(m_add[22]), .b(N134), .c(m_sub[22]), .d(N137), .out(n95) );
  aoi22 U173 ( .a(m_mul[22]), .b(N140), .c(m_kro[22]), .d(n14), .out(n94) );
  nand2 U174 ( .a(n96), .b(n97), .out(N26) );
  aoi22 U175 ( .a(m_add[21]), .b(N134), .c(m_sub[21]), .d(N137), .out(n97) );
  aoi22 U176 ( .a(m_mul[21]), .b(N140), .c(m_kro[21]), .d(n14), .out(n96) );
  nand2 U177 ( .a(n98), .b(n99), .out(N25) );
  aoi22 U178 ( .a(m_add[20]), .b(N134), .c(m_sub[20]), .d(N137), .out(n99) );
  aoi22 U179 ( .a(m_mul[20]), .b(N140), .c(m_kro[20]), .d(n14), .out(n98) );
  nand2 U180 ( .a(n100), .b(n101), .out(N24) );
  aoi22 U181 ( .a(m_add[19]), .b(N134), .c(m_sub[19]), .d(N137), .out(n101) );
  aoi22 U182 ( .a(m_mul[19]), .b(N140), .c(m_kro[19]), .d(n14), .out(n100) );
  nand2 U183 ( .a(n102), .b(n103), .out(N23) );
  aoi22 U184 ( .a(m_add[18]), .b(N134), .c(m_sub[18]), .d(N137), .out(n103) );
  aoi22 U185 ( .a(m_mul[18]), .b(N140), .c(m_kro[18]), .d(n14), .out(n102) );
  nand2 U186 ( .a(n104), .b(n105), .out(N22) );
  aoi22 U187 ( .a(m_add[17]), .b(N134), .c(m_sub[17]), .d(N137), .out(n105) );
  aoi22 U188 ( .a(m_mul[17]), .b(N140), .c(m_kro[17]), .d(n14), .out(n104) );
  nand2 U189 ( .a(n106), .b(n107), .out(N21) );
  aoi22 U190 ( .a(m_add[16]), .b(N134), .c(m_sub[16]), .d(N137), .out(n107) );
  aoi22 U191 ( .a(m_mul[16]), .b(N140), .c(m_kro[16]), .d(n14), .out(n106) );
  nand2 U192 ( .a(n108), .b(n109), .out(N20) );
  aoi22 U193 ( .a(m_add[15]), .b(N134), .c(m_sub[15]), .d(N137), .out(n109) );
  aoi22 U194 ( .a(m_mul[15]), .b(N140), .c(m_kro[15]), .d(n14), .out(n108) );
  nand2 U195 ( .a(n110), .b(n111), .out(N19) );
  aoi22 U196 ( .a(m_add[14]), .b(N134), .c(m_sub[14]), .d(N137), .out(n111) );
  aoi22 U197 ( .a(m_mul[14]), .b(N140), .c(m_kro[14]), .d(n14), .out(n110) );
  nand2 U198 ( .a(n112), .b(n113), .out(N18) );
  aoi22 U199 ( .a(m_add[13]), .b(N134), .c(m_sub[13]), .d(N137), .out(n113) );
  aoi22 U200 ( .a(m_mul[13]), .b(N140), .c(m_kro[13]), .d(n14), .out(n112) );
  nand2 U201 ( .a(n114), .b(n115), .out(N17) );
  aoi22 U202 ( .a(m_add[12]), .b(N134), .c(m_sub[12]), .d(N137), .out(n115) );
  aoi22 U203 ( .a(m_mul[12]), .b(N140), .c(m_kro[12]), .d(n14), .out(n114) );
  nand2 U204 ( .a(n116), .b(n117), .out(N16) );
  aoi22 U205 ( .a(m_add[11]), .b(N134), .c(m_sub[11]), .d(N137), .out(n117) );
  aoi22 U206 ( .a(m_mul[11]), .b(N140), .c(m_kro[11]), .d(n14), .out(n116) );
  nand2 U207 ( .a(n118), .b(n119), .out(N15) );
  aoi22 U208 ( .a(m_add[10]), .b(N134), .c(m_sub[10]), .d(N137), .out(n119) );
  aoi22 U209 ( .a(m_mul[10]), .b(N140), .c(m_kro[10]), .d(n14), .out(n118) );
  nand2 U210 ( .a(n120), .b(n121), .out(N14) );
  aoi22 U211 ( .a(m_add[9]), .b(N134), .c(m_sub[9]), .d(N137), .out(n121) );
  aoi22 U212 ( .a(m_mul[9]), .b(N140), .c(m_kro[9]), .d(n14), .out(n120) );
  nor2 U213 ( .a(n1), .b(n122), .out(N132) );
  inv U214 ( .in(m_kro[127]), .out(n122) );
  nor2 U215 ( .a(n1), .b(n123), .out(N131) );
  inv U216 ( .in(m_kro[126]), .out(n123) );
  nor2 U217 ( .a(n1), .b(n124), .out(N130) );
  inv U218 ( .in(m_kro[125]), .out(n124) );
  nand2 U219 ( .a(n125), .b(n126), .out(N13) );
  aoi22 U220 ( .a(m_add[8]), .b(N134), .c(m_sub[8]), .d(N137), .out(n126) );
  aoi22 U221 ( .a(m_mul[8]), .b(N140), .c(m_kro[8]), .d(n14), .out(n125) );
  nor2 U222 ( .a(n1), .b(n127), .out(N129) );
  inv U223 ( .in(m_kro[124]), .out(n127) );
  nor2 U224 ( .a(n1), .b(n128), .out(N128) );
  inv U225 ( .in(m_kro[123]), .out(n128) );
  nor2 U226 ( .a(n1), .b(n129), .out(N127) );
  inv U227 ( .in(m_kro[122]), .out(n129) );
  nor2 U228 ( .a(n1), .b(n130), .out(N126) );
  inv U229 ( .in(m_kro[121]), .out(n130) );
  nor2 U230 ( .a(n1), .b(n131), .out(N125) );
  inv U231 ( .in(m_kro[120]), .out(n131) );
  nor2 U232 ( .a(n1), .b(n132), .out(N124) );
  inv U233 ( .in(m_kro[119]), .out(n132) );
  nor2 U234 ( .a(n1), .b(n133), .out(N123) );
  inv U235 ( .in(m_kro[118]), .out(n133) );
  nor2 U236 ( .a(n1), .b(n134), .out(N122) );
  inv U237 ( .in(m_kro[117]), .out(n134) );
  nor2 U238 ( .a(n1), .b(n135), .out(N121) );
  inv U239 ( .in(m_kro[116]), .out(n135) );
  nor2 U240 ( .a(n1), .b(n136), .out(N120) );
  inv U241 ( .in(m_kro[115]), .out(n136) );
  nand2 U242 ( .a(n137), .b(n138), .out(N12) );
  aoi22 U243 ( .a(m_add[7]), .b(N134), .c(m_sub[7]), .d(N137), .out(n138) );
  aoi22 U244 ( .a(m_mul[7]), .b(N140), .c(m_kro[7]), .d(n14), .out(n137) );
  nor2 U245 ( .a(n1), .b(n139), .out(N119) );
  inv U246 ( .in(m_kro[114]), .out(n139) );
  nor2 U247 ( .a(n1), .b(n140), .out(N118) );
  inv U248 ( .in(m_kro[113]), .out(n140) );
  nor2 U249 ( .a(n1), .b(n141), .out(N117) );
  inv U250 ( .in(m_kro[112]), .out(n141) );
  nor2 U251 ( .a(n1), .b(n142), .out(N116) );
  inv U252 ( .in(m_kro[111]), .out(n142) );
  nor2 U253 ( .a(n1), .b(n143), .out(N115) );
  inv U254 ( .in(m_kro[110]), .out(n143) );
  nor2 U255 ( .a(n1), .b(n144), .out(N114) );
  inv U256 ( .in(m_kro[109]), .out(n144) );
  nor2 U257 ( .a(n1), .b(n145), .out(N113) );
  inv U258 ( .in(m_kro[108]), .out(n145) );
  nor2 U259 ( .a(n1), .b(n146), .out(N112) );
  inv U260 ( .in(m_kro[107]), .out(n146) );
  nor2 U261 ( .a(n1), .b(n147), .out(N111) );
  inv U262 ( .in(m_kro[106]), .out(n147) );
  nor2 U263 ( .a(n1), .b(n148), .out(N110) );
  inv U264 ( .in(m_kro[105]), .out(n148) );
  nand2 U265 ( .a(n149), .b(n150), .out(N11) );
  aoi22 U266 ( .a(m_add[6]), .b(N134), .c(m_sub[6]), .d(N137), .out(n150) );
  aoi22 U267 ( .a(m_mul[6]), .b(N140), .c(m_kro[6]), .d(n14), .out(n149) );
  nor2 U268 ( .a(n1), .b(n151), .out(N109) );
  inv U269 ( .in(m_kro[104]), .out(n151) );
  nor2 U270 ( .a(n1), .b(n152), .out(N108) );
  inv U271 ( .in(m_kro[103]), .out(n152) );
  nor2 U272 ( .a(n1), .b(n153), .out(N107) );
  inv U273 ( .in(m_kro[102]), .out(n153) );
  nor2 U274 ( .a(n1), .b(n154), .out(N106) );
  inv U275 ( .in(m_kro[101]), .out(n154) );
  nor2 U276 ( .a(n1), .b(n155), .out(N105) );
  inv U277 ( .in(m_kro[100]), .out(n155) );
  nor2 U278 ( .a(n1), .b(n156), .out(N104) );
  inv U279 ( .in(m_kro[99]), .out(n156) );
  nor2 U280 ( .a(n1), .b(n157), .out(N103) );
  inv U281 ( .in(m_kro[98]), .out(n157) );
  nor2 U282 ( .a(n1), .b(n158), .out(N102) );
  inv U283 ( .in(m_kro[97]), .out(n158) );
  nor2 U284 ( .a(n1), .b(n159), .out(N101) );
  inv U285 ( .in(m_kro[96]), .out(n159) );
  nor2 U286 ( .a(n1), .b(n160), .out(N100) );
  inv U287 ( .in(m_kro[95]), .out(n160) );
  nand2 U288 ( .a(n161), .b(n162), .out(N10) );
  aoi22 U289 ( .a(m_add[5]), .b(N134), .c(m_sub[5]), .d(N137), .out(n162) );
  aoi22 U290 ( .a(m_mul[5]), .b(N140), .c(m_kro[5]), .d(n14), .out(n161) );
  inv U291 ( .in(n1), .out(n14) );
  inv U292 ( .in(op[1]), .out(n163) );
  inv \mat_kron/mult_40/AN1_7  ( .in(A[31]), .out(\mat_kron/mult_40/A_not [7])
         );
  inv \mat_kron/mult_40/AN1_6  ( .in(A[30]), .out(\mat_kron/mult_40/A_not [6])
         );
  inv \mat_kron/mult_40/AN1_5  ( .in(A[29]), .out(\mat_kron/mult_40/A_not [5])
         );
  inv \mat_kron/mult_40/AN1_4  ( .in(A[28]), .out(\mat_kron/mult_40/A_not [4])
         );
  inv \mat_kron/mult_40/AN1_3  ( .in(A[27]), .out(\mat_kron/mult_40/A_not [3])
         );
  inv \mat_kron/mult_40/AN1_2  ( .in(A[26]), .out(\mat_kron/mult_40/A_not [2])
         );
  inv \mat_kron/mult_40/AN1_1  ( .in(A[25]), .out(\mat_kron/mult_40/A_not [1])
         );
  inv \mat_kron/mult_40/AN1_0  ( .in(A[24]), .out(\mat_kron/mult_40/A_notx[0] ) );
  inv \mat_kron/mult_40/AN1_7_0  ( .in(\mat_add/r94/B_AS [7]), .out(
        \mat_kron/mult_40/B_not [7]) );
  inv \mat_kron/mult_40/AN1_6_0  ( .in(\mat_add/r94/B_AS [6]), .out(
        \mat_kron/mult_40/B_not [6]) );
  inv \mat_kron/mult_40/AN1_5_0  ( .in(\mat_add/r94/B_AS [5]), .out(
        \mat_kron/mult_40/B_not [5]) );
  inv \mat_kron/mult_40/AN1_4_0  ( .in(\mat_add/r94/B_AS [4]), .out(
        \mat_kron/mult_40/B_not [4]) );
  inv \mat_kron/mult_40/AN1_3_0  ( .in(\mat_add/r94/B_AS [3]), .out(
        \mat_kron/mult_40/B_not [3]) );
  inv \mat_kron/mult_40/AN1_2_0  ( .in(\mat_add/r94/B_AS [2]), .out(
        \mat_kron/mult_40/B_not [2]) );
  inv \mat_kron/mult_40/AN1_1_0  ( .in(\mat_add/r94/B_AS [1]), .out(
        \mat_kron/mult_40/B_not [1]) );
  inv \mat_kron/mult_40/AN1_0_0  ( .in(\mat_add/r94/B_AS [0]), .out(
        \mat_kron/mult_40/B_notx[0] ) );
  nor2 \mat_kron/mult_40/AN3_7_0  ( .a(\mat_kron/mult_40/A_not [7]), .b(
        \mat_kron/mult_40/B_notx[0] ), .out(\mat_kron/mult_40/ab[7][0] ) );
  nor2 \mat_kron/mult_40/AN1_6_1  ( .a(\mat_kron/mult_40/A_not [6]), .b(
        \mat_kron/mult_40/B_not [1]), .out(\mat_kron/mult_40/ab[6][1] ) );
  nor2 \mat_kron/mult_40/AN1_6_0_0  ( .a(\mat_kron/mult_40/A_not [6]), .b(
        \mat_kron/mult_40/B_notx[0] ), .out(\mat_kron/mult_40/ab[6][0] ) );
  nor2 \mat_kron/mult_40/AN1_5_2  ( .a(\mat_kron/mult_40/A_not [5]), .b(
        \mat_kron/mult_40/B_not [2]), .out(\mat_kron/mult_40/ab[5][2] ) );
  nor2 \mat_kron/mult_40/AN1_5_1  ( .a(\mat_kron/mult_40/A_not [5]), .b(
        \mat_kron/mult_40/B_not [1]), .out(\mat_kron/mult_40/ab[5][1] ) );
  nor2 \mat_kron/mult_40/AN1_5_0_0  ( .a(\mat_kron/mult_40/A_not [5]), .b(
        \mat_kron/mult_40/B_notx[0] ), .out(\mat_kron/mult_40/ab[5][0] ) );
  nor2 \mat_kron/mult_40/AN1_4_3  ( .a(\mat_kron/mult_40/A_not [4]), .b(
        \mat_kron/mult_40/B_not [3]), .out(\mat_kron/mult_40/ab[4][3] ) );
  nor2 \mat_kron/mult_40/AN1_4_2  ( .a(\mat_kron/mult_40/A_not [4]), .b(
        \mat_kron/mult_40/B_not [2]), .out(\mat_kron/mult_40/ab[4][2] ) );
  nor2 \mat_kron/mult_40/AN1_4_1  ( .a(\mat_kron/mult_40/A_not [4]), .b(
        \mat_kron/mult_40/B_not [1]), .out(\mat_kron/mult_40/ab[4][1] ) );
  nor2 \mat_kron/mult_40/AN1_4_0_0  ( .a(\mat_kron/mult_40/A_not [4]), .b(
        \mat_kron/mult_40/B_notx[0] ), .out(\mat_kron/mult_40/ab[4][0] ) );
  nor2 \mat_kron/mult_40/AN1_3_4  ( .a(\mat_kron/mult_40/A_not [3]), .b(
        \mat_kron/mult_40/B_not [4]), .out(\mat_kron/mult_40/ab[3][4] ) );
  nor2 \mat_kron/mult_40/AN1_3_3  ( .a(\mat_kron/mult_40/A_not [3]), .b(
        \mat_kron/mult_40/B_not [3]), .out(\mat_kron/mult_40/ab[3][3] ) );
  nor2 \mat_kron/mult_40/AN1_3_2  ( .a(\mat_kron/mult_40/A_not [3]), .b(
        \mat_kron/mult_40/B_not [2]), .out(\mat_kron/mult_40/ab[3][2] ) );
  nor2 \mat_kron/mult_40/AN1_3_1  ( .a(\mat_kron/mult_40/A_not [3]), .b(
        \mat_kron/mult_40/B_not [1]), .out(\mat_kron/mult_40/ab[3][1] ) );
  nor2 \mat_kron/mult_40/AN1_3_0_0  ( .a(\mat_kron/mult_40/A_not [3]), .b(
        \mat_kron/mult_40/B_notx[0] ), .out(\mat_kron/mult_40/ab[3][0] ) );
  nor2 \mat_kron/mult_40/AN1_2_5  ( .a(\mat_kron/mult_40/A_not [2]), .b(
        \mat_kron/mult_40/B_not [5]), .out(\mat_kron/mult_40/ab[2][5] ) );
  nor2 \mat_kron/mult_40/AN1_2_4  ( .a(\mat_kron/mult_40/A_not [2]), .b(
        \mat_kron/mult_40/B_not [4]), .out(\mat_kron/mult_40/ab[2][4] ) );
  nor2 \mat_kron/mult_40/AN1_2_3  ( .a(\mat_kron/mult_40/A_not [2]), .b(
        \mat_kron/mult_40/B_not [3]), .out(\mat_kron/mult_40/ab[2][3] ) );
  nor2 \mat_kron/mult_40/AN1_2_2  ( .a(\mat_kron/mult_40/A_not [2]), .b(
        \mat_kron/mult_40/B_not [2]), .out(\mat_kron/mult_40/ab[2][2] ) );
  nor2 \mat_kron/mult_40/AN1_2_1  ( .a(\mat_kron/mult_40/A_not [2]), .b(
        \mat_kron/mult_40/B_not [1]), .out(\mat_kron/mult_40/ab[2][1] ) );
  nor2 \mat_kron/mult_40/AN1_2_0_0  ( .a(\mat_kron/mult_40/A_not [2]), .b(
        \mat_kron/mult_40/B_notx[0] ), .out(\mat_kron/mult_40/ab[2][0] ) );
  nor2 \mat_kron/mult_40/AN1_1_6  ( .a(\mat_kron/mult_40/A_not [1]), .b(
        \mat_kron/mult_40/B_not [6]), .out(\mat_kron/mult_40/ab[1][6] ) );
  nor2 \mat_kron/mult_40/AN1_1_5  ( .a(\mat_kron/mult_40/A_not [1]), .b(
        \mat_kron/mult_40/B_not [5]), .out(\mat_kron/mult_40/ab[1][5] ) );
  nor2 \mat_kron/mult_40/AN1_1_4  ( .a(\mat_kron/mult_40/A_not [1]), .b(
        \mat_kron/mult_40/B_not [4]), .out(\mat_kron/mult_40/ab[1][4] ) );
  nor2 \mat_kron/mult_40/AN1_1_3  ( .a(\mat_kron/mult_40/A_not [1]), .b(
        \mat_kron/mult_40/B_not [3]), .out(\mat_kron/mult_40/ab[1][3] ) );
  nor2 \mat_kron/mult_40/AN1_1_2  ( .a(\mat_kron/mult_40/A_not [1]), .b(
        \mat_kron/mult_40/B_not [2]), .out(\mat_kron/mult_40/ab[1][2] ) );
  nor2 \mat_kron/mult_40/AN1_1_1  ( .a(\mat_kron/mult_40/A_not [1]), .b(
        \mat_kron/mult_40/B_not [1]), .out(\mat_kron/mult_40/ab[1][1] ) );
  nor2 \mat_kron/mult_40/AN1_1_0_0  ( .a(\mat_kron/mult_40/A_not [1]), .b(
        \mat_kron/mult_40/B_notx[0] ), .out(\mat_kron/mult_40/ab[1][0] ) );
  nor2 \mat_kron/mult_40/AN2_0_7  ( .a(\mat_kron/mult_40/A_notx[0] ), .b(
        \mat_kron/mult_40/B_not [7]), .out(\mat_kron/mult_40/ab[0][7] ) );
  nor2 \mat_kron/mult_40/AN1_0_6  ( .a(\mat_kron/mult_40/A_notx[0] ), .b(
        \mat_kron/mult_40/B_not [6]), .out(\mat_kron/mult_40/ab[0][6] ) );
  nor2 \mat_kron/mult_40/AN1_0_5  ( .a(\mat_kron/mult_40/A_notx[0] ), .b(
        \mat_kron/mult_40/B_not [5]), .out(\mat_kron/mult_40/ab[0][5] ) );
  nor2 \mat_kron/mult_40/AN1_0_4  ( .a(\mat_kron/mult_40/A_notx[0] ), .b(
        \mat_kron/mult_40/B_not [4]), .out(\mat_kron/mult_40/ab[0][4] ) );
  nor2 \mat_kron/mult_40/AN1_0_3  ( .a(\mat_kron/mult_40/A_notx[0] ), .b(
        \mat_kron/mult_40/B_not [3]), .out(\mat_kron/mult_40/ab[0][3] ) );
  nor2 \mat_kron/mult_40/AN1_0_2  ( .a(\mat_kron/mult_40/A_notx[0] ), .b(
        \mat_kron/mult_40/B_not [2]), .out(\mat_kron/mult_40/ab[0][2] ) );
  nor2 \mat_kron/mult_40/AN1_0_1  ( .a(\mat_kron/mult_40/A_notx[0] ), .b(
        \mat_kron/mult_40/B_not [1]), .out(\mat_kron/mult_40/ab[0][1] ) );
  nor2 \mat_kron/mult_40/AN1_0_0_0  ( .a(\mat_kron/mult_40/A_notx[0] ), .b(
        \mat_kron/mult_40/B_notx[0] ), .out(m_kro[120]) );
  inv \mat_kron/mult_40_G2_G1_G1_G1/AN1_7  ( .in(A[31]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [7]) );
  inv \mat_kron/mult_40_G2_G1_G1_G1/AN1_6  ( .in(A[30]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [6]) );
  inv \mat_kron/mult_40_G2_G1_G1_G1/AN1_5  ( .in(A[29]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [5]) );
  inv \mat_kron/mult_40_G2_G1_G1_G1/AN1_4  ( .in(A[28]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [4]) );
  inv \mat_kron/mult_40_G2_G1_G1_G1/AN1_3  ( .in(A[27]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [3]) );
  inv \mat_kron/mult_40_G2_G1_G1_G1/AN1_2  ( .in(A[26]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [2]) );
  inv \mat_kron/mult_40_G2_G1_G1_G1/AN1_1  ( .in(A[25]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [1]) );
  inv \mat_kron/mult_40_G2_G1_G1_G1/AN1_0  ( .in(A[24]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/A_notx[0] ) );
  inv \mat_kron/mult_40_G2_G1_G1_G1/AN1_7_0  ( .in(\mat_add/r98/B_AS [7]), 
        .out(\mat_kron/mult_40_G2_G1_G1_G1/B_not [7]) );
  inv \mat_kron/mult_40_G2_G1_G1_G1/AN1_6_0  ( .in(\mat_add/r98/B_AS [6]), 
        .out(\mat_kron/mult_40_G2_G1_G1_G1/B_not [6]) );
  inv \mat_kron/mult_40_G2_G1_G1_G1/AN1_5_0  ( .in(\mat_add/r98/B_AS [5]), 
        .out(\mat_kron/mult_40_G2_G1_G1_G1/B_not [5]) );
  inv \mat_kron/mult_40_G2_G1_G1_G1/AN1_4_0  ( .in(\mat_add/r98/B_AS [4]), 
        .out(\mat_kron/mult_40_G2_G1_G1_G1/B_not [4]) );
  inv \mat_kron/mult_40_G2_G1_G1_G1/AN1_3_0  ( .in(\mat_add/r98/B_AS [3]), 
        .out(\mat_kron/mult_40_G2_G1_G1_G1/B_not [3]) );
  inv \mat_kron/mult_40_G2_G1_G1_G1/AN1_2_0  ( .in(\mat_add/r98/B_AS [2]), 
        .out(\mat_kron/mult_40_G2_G1_G1_G1/B_not [2]) );
  inv \mat_kron/mult_40_G2_G1_G1_G1/AN1_1_0  ( .in(\mat_add/r98/B_AS [1]), 
        .out(\mat_kron/mult_40_G2_G1_G1_G1/B_not [1]) );
  inv \mat_kron/mult_40_G2_G1_G1_G1/AN1_0_0  ( .in(\mat_add/r98/B_AS [0]), 
        .out(\mat_kron/mult_40_G2_G1_G1_G1/B_notx[0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN3_7_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [7]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[7][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_6_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [6]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[6][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_6_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [6]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[6][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_5_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[5][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_5_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[5][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_5_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[5][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_4_3  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[4][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_4_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[4][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_4_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[4][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_4_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[4][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_3_4  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[3][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_3_3  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[3][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_3_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[3][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_3_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[3][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_3_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[3][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_2_5  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[2][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_2_4  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[2][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_2_3  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[2][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_2_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[2][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_2_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[2][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_2_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[2][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_1_6  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [6]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[1][6] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_1_5  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[1][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_1_4  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[1][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_1_3  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[1][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_1_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[1][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_1_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[1][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_1_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[1][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN2_0_7  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [7]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[0][7] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_0_6  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [6]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[0][6] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_0_5  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[0][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_0_4  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[0][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_0_3  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[0][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_0_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[0][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_0_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[0][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G1/AN1_0_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/B_notx[0] ), .out(m_kro[112]) );
  inv \mat_kron/mult_40_G2_G1_G1/AN1_7  ( .in(A[31]), .out(
        \mat_kron/mult_40_G2_G1_G1/A_not [7]) );
  inv \mat_kron/mult_40_G2_G1_G1/AN1_6  ( .in(A[30]), .out(
        \mat_kron/mult_40_G2_G1_G1/A_not [6]) );
  inv \mat_kron/mult_40_G2_G1_G1/AN1_5  ( .in(A[29]), .out(
        \mat_kron/mult_40_G2_G1_G1/A_not [5]) );
  inv \mat_kron/mult_40_G2_G1_G1/AN1_4  ( .in(A[28]), .out(
        \mat_kron/mult_40_G2_G1_G1/A_not [4]) );
  inv \mat_kron/mult_40_G2_G1_G1/AN1_3  ( .in(A[27]), .out(
        \mat_kron/mult_40_G2_G1_G1/A_not [3]) );
  inv \mat_kron/mult_40_G2_G1_G1/AN1_2  ( .in(A[26]), .out(
        \mat_kron/mult_40_G2_G1_G1/A_not [2]) );
  inv \mat_kron/mult_40_G2_G1_G1/AN1_1  ( .in(A[25]), .out(
        \mat_kron/mult_40_G2_G1_G1/A_not [1]) );
  inv \mat_kron/mult_40_G2_G1_G1/AN1_0  ( .in(A[24]), .out(
        \mat_kron/mult_40_G2_G1_G1/A_notx[0] ) );
  inv \mat_kron/mult_40_G2_G1_G1/AN1_7_0  ( .in(\mat_add/r102/B_AS [7]), .out(
        \mat_kron/mult_40_G2_G1_G1/B_not [7]) );
  inv \mat_kron/mult_40_G2_G1_G1/AN1_6_0  ( .in(\mat_add/r102/B_AS [6]), .out(
        \mat_kron/mult_40_G2_G1_G1/B_not [6]) );
  inv \mat_kron/mult_40_G2_G1_G1/AN1_5_0  ( .in(\mat_add/r102/B_AS [5]), .out(
        \mat_kron/mult_40_G2_G1_G1/B_not [5]) );
  inv \mat_kron/mult_40_G2_G1_G1/AN1_4_0  ( .in(\mat_add/r102/B_AS [4]), .out(
        \mat_kron/mult_40_G2_G1_G1/B_not [4]) );
  inv \mat_kron/mult_40_G2_G1_G1/AN1_3_0  ( .in(\mat_add/r102/B_AS [3]), .out(
        \mat_kron/mult_40_G2_G1_G1/B_not [3]) );
  inv \mat_kron/mult_40_G2_G1_G1/AN1_2_0  ( .in(\mat_add/r102/B_AS [2]), .out(
        \mat_kron/mult_40_G2_G1_G1/B_not [2]) );
  inv \mat_kron/mult_40_G2_G1_G1/AN1_1_0  ( .in(\mat_add/r102/B_AS [1]), .out(
        \mat_kron/mult_40_G2_G1_G1/B_not [1]) );
  inv \mat_kron/mult_40_G2_G1_G1/AN1_0_0  ( .in(\mat_add/r102/B_AS [0]), .out(
        \mat_kron/mult_40_G2_G1_G1/B_notx[0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN3_7_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [7]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[7][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_6_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [6]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[6][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_6_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [6]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[6][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_5_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[5][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_5_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[5][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_5_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[5][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_4_3  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[4][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_4_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[4][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_4_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[4][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_4_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[4][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_3_4  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[3][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_3_3  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[3][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_3_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[3][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_3_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[3][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_3_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[3][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_2_5  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[2][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_2_4  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[2][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_2_3  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[2][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_2_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[2][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_2_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[2][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_2_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[2][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_1_6  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [6]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[1][6] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_1_5  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[1][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_1_4  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[1][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_1_3  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[1][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_1_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[1][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_1_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[1][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_1_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[1][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN2_0_7  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [7]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[0][7] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_0_6  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [6]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[0][6] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_0_5  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[0][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_0_4  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[0][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_0_3  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[0][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_0_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[0][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_0_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1/ab[0][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1/AN1_0_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1/B_notx[0] ), .out(m_kro[88]) );
  inv \mat_kron/mult_40_G2_G2_G1_G1/AN1_7  ( .in(A[31]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [7]) );
  inv \mat_kron/mult_40_G2_G2_G1_G1/AN1_6  ( .in(A[30]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [6]) );
  inv \mat_kron/mult_40_G2_G2_G1_G1/AN1_5  ( .in(A[29]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [5]) );
  inv \mat_kron/mult_40_G2_G2_G1_G1/AN1_4  ( .in(A[28]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [4]) );
  inv \mat_kron/mult_40_G2_G2_G1_G1/AN1_3  ( .in(A[27]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [3]) );
  inv \mat_kron/mult_40_G2_G2_G1_G1/AN1_2  ( .in(A[26]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [2]) );
  inv \mat_kron/mult_40_G2_G2_G1_G1/AN1_1  ( .in(A[25]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [1]) );
  inv \mat_kron/mult_40_G2_G2_G1_G1/AN1_0  ( .in(A[24]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/A_notx[0] ) );
  inv \mat_kron/mult_40_G2_G2_G1_G1/AN1_7_0  ( .in(\mat_add/r106/B_AS [7]), 
        .out(\mat_kron/mult_40_G2_G2_G1_G1/B_not [7]) );
  inv \mat_kron/mult_40_G2_G2_G1_G1/AN1_6_0  ( .in(\mat_add/r106/B_AS [6]), 
        .out(\mat_kron/mult_40_G2_G2_G1_G1/B_not [6]) );
  inv \mat_kron/mult_40_G2_G2_G1_G1/AN1_5_0  ( .in(\mat_add/r106/B_AS [5]), 
        .out(\mat_kron/mult_40_G2_G2_G1_G1/B_not [5]) );
  inv \mat_kron/mult_40_G2_G2_G1_G1/AN1_4_0  ( .in(\mat_add/r106/B_AS [4]), 
        .out(\mat_kron/mult_40_G2_G2_G1_G1/B_not [4]) );
  inv \mat_kron/mult_40_G2_G2_G1_G1/AN1_3_0  ( .in(\mat_add/r106/B_AS [3]), 
        .out(\mat_kron/mult_40_G2_G2_G1_G1/B_not [3]) );
  inv \mat_kron/mult_40_G2_G2_G1_G1/AN1_2_0  ( .in(\mat_add/r106/B_AS [2]), 
        .out(\mat_kron/mult_40_G2_G2_G1_G1/B_not [2]) );
  inv \mat_kron/mult_40_G2_G2_G1_G1/AN1_1_0  ( .in(\mat_add/r106/B_AS [1]), 
        .out(\mat_kron/mult_40_G2_G2_G1_G1/B_not [1]) );
  inv \mat_kron/mult_40_G2_G2_G1_G1/AN1_0_0  ( .in(\mat_add/r106/B_AS [0]), 
        .out(\mat_kron/mult_40_G2_G2_G1_G1/B_notx[0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN3_7_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [7]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[7][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_6_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [6]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[6][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_6_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [6]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[6][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_5_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[5][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_5_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[5][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_5_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[5][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_4_3  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[4][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_4_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[4][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_4_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[4][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_4_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[4][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_3_4  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[3][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_3_3  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[3][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_3_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[3][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_3_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[3][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_3_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[3][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_2_5  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[2][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_2_4  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[2][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_2_3  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[2][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_2_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[2][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_2_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[2][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_2_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[2][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_1_6  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [6]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[1][6] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_1_5  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[1][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_1_4  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[1][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_1_3  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[1][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_1_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[1][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_1_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[1][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_1_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[1][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN2_0_7  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [7]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[0][7] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_0_6  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [6]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[0][6] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_0_5  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[0][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_0_4  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[0][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_0_3  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[0][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_0_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[0][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_0_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[0][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G1/AN1_0_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/B_notx[0] ), .out(m_kro[80]) );
  inv \mat_kron/mult_40_G2_G1/AN1_7  ( .in(A[23]), .out(
        \mat_kron/mult_40_G2_G1/A_not [7]) );
  inv \mat_kron/mult_40_G2_G1/AN1_6  ( .in(A[22]), .out(
        \mat_kron/mult_40_G2_G1/A_not [6]) );
  inv \mat_kron/mult_40_G2_G1/AN1_5  ( .in(A[21]), .out(
        \mat_kron/mult_40_G2_G1/A_not [5]) );
  inv \mat_kron/mult_40_G2_G1/AN1_4  ( .in(A[20]), .out(
        \mat_kron/mult_40_G2_G1/A_not [4]) );
  inv \mat_kron/mult_40_G2_G1/AN1_3  ( .in(A[19]), .out(
        \mat_kron/mult_40_G2_G1/A_not [3]) );
  inv \mat_kron/mult_40_G2_G1/AN1_2  ( .in(A[18]), .out(
        \mat_kron/mult_40_G2_G1/A_not [2]) );
  inv \mat_kron/mult_40_G2_G1/AN1_1  ( .in(A[17]), .out(
        \mat_kron/mult_40_G2_G1/A_not [1]) );
  inv \mat_kron/mult_40_G2_G1/AN1_0  ( .in(A[16]), .out(
        \mat_kron/mult_40_G2_G1/A_notx[0] ) );
  inv \mat_kron/mult_40_G2_G1/AN1_7_0  ( .in(\mat_add/r94/B_AS [7]), .out(
        \mat_kron/mult_40_G2_G1/B_not [7]) );
  inv \mat_kron/mult_40_G2_G1/AN1_6_0  ( .in(\mat_add/r94/B_AS [6]), .out(
        \mat_kron/mult_40_G2_G1/B_not [6]) );
  inv \mat_kron/mult_40_G2_G1/AN1_5_0  ( .in(\mat_add/r94/B_AS [5]), .out(
        \mat_kron/mult_40_G2_G1/B_not [5]) );
  inv \mat_kron/mult_40_G2_G1/AN1_4_0  ( .in(\mat_add/r94/B_AS [4]), .out(
        \mat_kron/mult_40_G2_G1/B_not [4]) );
  inv \mat_kron/mult_40_G2_G1/AN1_3_0  ( .in(\mat_add/r94/B_AS [3]), .out(
        \mat_kron/mult_40_G2_G1/B_not [3]) );
  inv \mat_kron/mult_40_G2_G1/AN1_2_0  ( .in(\mat_add/r94/B_AS [2]), .out(
        \mat_kron/mult_40_G2_G1/B_not [2]) );
  inv \mat_kron/mult_40_G2_G1/AN1_1_0  ( .in(\mat_add/r94/B_AS [1]), .out(
        \mat_kron/mult_40_G2_G1/B_not [1]) );
  inv \mat_kron/mult_40_G2_G1/AN1_0_0  ( .in(\mat_add/r94/B_AS [0]), .out(
        \mat_kron/mult_40_G2_G1/B_notx[0] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN3_7_0  ( .a(\mat_kron/mult_40_G2_G1/A_not [7]), .b(\mat_kron/mult_40_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1/ab[7][0] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_6_1  ( .a(\mat_kron/mult_40_G2_G1/A_not [6]), .b(\mat_kron/mult_40_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1/ab[6][1] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_6_0_0  ( .a(
        \mat_kron/mult_40_G2_G1/A_not [6]), .b(
        \mat_kron/mult_40_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1/ab[6][0] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_5_2  ( .a(\mat_kron/mult_40_G2_G1/A_not [5]), .b(\mat_kron/mult_40_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1/ab[5][2] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_5_1  ( .a(\mat_kron/mult_40_G2_G1/A_not [5]), .b(\mat_kron/mult_40_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1/ab[5][1] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_5_0_0  ( .a(
        \mat_kron/mult_40_G2_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1/ab[5][0] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_4_3  ( .a(\mat_kron/mult_40_G2_G1/A_not [4]), .b(\mat_kron/mult_40_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1/ab[4][3] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_4_2  ( .a(\mat_kron/mult_40_G2_G1/A_not [4]), .b(\mat_kron/mult_40_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1/ab[4][2] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_4_1  ( .a(\mat_kron/mult_40_G2_G1/A_not [4]), .b(\mat_kron/mult_40_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1/ab[4][1] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_4_0_0  ( .a(
        \mat_kron/mult_40_G2_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1/ab[4][0] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_3_4  ( .a(\mat_kron/mult_40_G2_G1/A_not [3]), .b(\mat_kron/mult_40_G2_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1/ab[3][4] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_3_3  ( .a(\mat_kron/mult_40_G2_G1/A_not [3]), .b(\mat_kron/mult_40_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1/ab[3][3] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_3_2  ( .a(\mat_kron/mult_40_G2_G1/A_not [3]), .b(\mat_kron/mult_40_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1/ab[3][2] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_3_1  ( .a(\mat_kron/mult_40_G2_G1/A_not [3]), .b(\mat_kron/mult_40_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1/ab[3][1] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_3_0_0  ( .a(
        \mat_kron/mult_40_G2_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1/ab[3][0] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_2_5  ( .a(\mat_kron/mult_40_G2_G1/A_not [2]), .b(\mat_kron/mult_40_G2_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1/ab[2][5] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_2_4  ( .a(\mat_kron/mult_40_G2_G1/A_not [2]), .b(\mat_kron/mult_40_G2_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1/ab[2][4] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_2_3  ( .a(\mat_kron/mult_40_G2_G1/A_not [2]), .b(\mat_kron/mult_40_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1/ab[2][3] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_2_2  ( .a(\mat_kron/mult_40_G2_G1/A_not [2]), .b(\mat_kron/mult_40_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1/ab[2][2] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_2_1  ( .a(\mat_kron/mult_40_G2_G1/A_not [2]), .b(\mat_kron/mult_40_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1/ab[2][1] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_2_0_0  ( .a(
        \mat_kron/mult_40_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1/ab[2][0] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_1_6  ( .a(\mat_kron/mult_40_G2_G1/A_not [1]), .b(\mat_kron/mult_40_G2_G1/B_not [6]), .out(
        \mat_kron/mult_40_G2_G1/ab[1][6] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_1_5  ( .a(\mat_kron/mult_40_G2_G1/A_not [1]), .b(\mat_kron/mult_40_G2_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1/ab[1][5] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_1_4  ( .a(\mat_kron/mult_40_G2_G1/A_not [1]), .b(\mat_kron/mult_40_G2_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1/ab[1][4] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_1_3  ( .a(\mat_kron/mult_40_G2_G1/A_not [1]), .b(\mat_kron/mult_40_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1/ab[1][3] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_1_2  ( .a(\mat_kron/mult_40_G2_G1/A_not [1]), .b(\mat_kron/mult_40_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1/ab[1][2] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_1_1  ( .a(\mat_kron/mult_40_G2_G1/A_not [1]), .b(\mat_kron/mult_40_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1/ab[1][1] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_1_0_0  ( .a(
        \mat_kron/mult_40_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1/ab[1][0] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN2_0_7  ( .a(
        \mat_kron/mult_40_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1/B_not [7]), .out(
        \mat_kron/mult_40_G2_G1/ab[0][7] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_0_6  ( .a(
        \mat_kron/mult_40_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1/B_not [6]), .out(
        \mat_kron/mult_40_G2_G1/ab[0][6] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_0_5  ( .a(
        \mat_kron/mult_40_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1/ab[0][5] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_0_4  ( .a(
        \mat_kron/mult_40_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1/ab[0][4] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_0_3  ( .a(
        \mat_kron/mult_40_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1/ab[0][3] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_0_2  ( .a(
        \mat_kron/mult_40_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1/ab[0][2] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_0_1  ( .a(
        \mat_kron/mult_40_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1/ab[0][1] ) );
  nor2 \mat_kron/mult_40_G2_G1/AN1_0_0_0  ( .a(
        \mat_kron/mult_40_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1/B_notx[0] ), .out(m_kro[104]) );
  inv \mat_kron/mult_40_G2_G1_G2_G1/AN1_7  ( .in(A[23]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [7]) );
  inv \mat_kron/mult_40_G2_G1_G2_G1/AN1_6  ( .in(A[22]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [6]) );
  inv \mat_kron/mult_40_G2_G1_G2_G1/AN1_5  ( .in(A[21]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [5]) );
  inv \mat_kron/mult_40_G2_G1_G2_G1/AN1_4  ( .in(A[20]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [4]) );
  inv \mat_kron/mult_40_G2_G1_G2_G1/AN1_3  ( .in(A[19]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [3]) );
  inv \mat_kron/mult_40_G2_G1_G2_G1/AN1_2  ( .in(A[18]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [2]) );
  inv \mat_kron/mult_40_G2_G1_G2_G1/AN1_1  ( .in(A[17]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [1]) );
  inv \mat_kron/mult_40_G2_G1_G2_G1/AN1_0  ( .in(A[16]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/A_notx[0] ) );
  inv \mat_kron/mult_40_G2_G1_G2_G1/AN1_7_0  ( .in(\mat_add/r98/B_AS [7]), 
        .out(\mat_kron/mult_40_G2_G1_G2_G1/B_not [7]) );
  inv \mat_kron/mult_40_G2_G1_G2_G1/AN1_6_0  ( .in(\mat_add/r98/B_AS [6]), 
        .out(\mat_kron/mult_40_G2_G1_G2_G1/B_not [6]) );
  inv \mat_kron/mult_40_G2_G1_G2_G1/AN1_5_0  ( .in(\mat_add/r98/B_AS [5]), 
        .out(\mat_kron/mult_40_G2_G1_G2_G1/B_not [5]) );
  inv \mat_kron/mult_40_G2_G1_G2_G1/AN1_4_0  ( .in(\mat_add/r98/B_AS [4]), 
        .out(\mat_kron/mult_40_G2_G1_G2_G1/B_not [4]) );
  inv \mat_kron/mult_40_G2_G1_G2_G1/AN1_3_0  ( .in(\mat_add/r98/B_AS [3]), 
        .out(\mat_kron/mult_40_G2_G1_G2_G1/B_not [3]) );
  inv \mat_kron/mult_40_G2_G1_G2_G1/AN1_2_0  ( .in(\mat_add/r98/B_AS [2]), 
        .out(\mat_kron/mult_40_G2_G1_G2_G1/B_not [2]) );
  inv \mat_kron/mult_40_G2_G1_G2_G1/AN1_1_0  ( .in(\mat_add/r98/B_AS [1]), 
        .out(\mat_kron/mult_40_G2_G1_G2_G1/B_not [1]) );
  inv \mat_kron/mult_40_G2_G1_G2_G1/AN1_0_0  ( .in(\mat_add/r98/B_AS [0]), 
        .out(\mat_kron/mult_40_G2_G1_G2_G1/B_notx[0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN3_7_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [7]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[7][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_6_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [6]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[6][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_6_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [6]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[6][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_5_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[5][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_5_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[5][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_5_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[5][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_4_3  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[4][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_4_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[4][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_4_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[4][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_4_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[4][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_3_4  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[3][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_3_3  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[3][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_3_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[3][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_3_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[3][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_3_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[3][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_2_5  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[2][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_2_4  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[2][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_2_3  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[2][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_2_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[2][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_2_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[2][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_2_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[2][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_1_6  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [6]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[1][6] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_1_5  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[1][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_1_4  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[1][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_1_3  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[1][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_1_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[1][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_1_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[1][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_1_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[1][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN2_0_7  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [7]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[0][7] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_0_6  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [6]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[0][6] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_0_5  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[0][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_0_4  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[0][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_0_3  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[0][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_0_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[0][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_0_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[0][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G1/AN1_0_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/B_notx[0] ), .out(m_kro[96]) );
  inv \mat_kron/mult_40_G2_G2_G1/AN1_7  ( .in(A[23]), .out(
        \mat_kron/mult_40_G2_G2_G1/A_not [7]) );
  inv \mat_kron/mult_40_G2_G2_G1/AN1_6  ( .in(A[22]), .out(
        \mat_kron/mult_40_G2_G2_G1/A_not [6]) );
  inv \mat_kron/mult_40_G2_G2_G1/AN1_5  ( .in(A[21]), .out(
        \mat_kron/mult_40_G2_G2_G1/A_not [5]) );
  inv \mat_kron/mult_40_G2_G2_G1/AN1_4  ( .in(A[20]), .out(
        \mat_kron/mult_40_G2_G2_G1/A_not [4]) );
  inv \mat_kron/mult_40_G2_G2_G1/AN1_3  ( .in(A[19]), .out(
        \mat_kron/mult_40_G2_G2_G1/A_not [3]) );
  inv \mat_kron/mult_40_G2_G2_G1/AN1_2  ( .in(A[18]), .out(
        \mat_kron/mult_40_G2_G2_G1/A_not [2]) );
  inv \mat_kron/mult_40_G2_G2_G1/AN1_1  ( .in(A[17]), .out(
        \mat_kron/mult_40_G2_G2_G1/A_not [1]) );
  inv \mat_kron/mult_40_G2_G2_G1/AN1_0  ( .in(A[16]), .out(
        \mat_kron/mult_40_G2_G2_G1/A_notx[0] ) );
  inv \mat_kron/mult_40_G2_G2_G1/AN1_7_0  ( .in(\mat_add/r102/B_AS [7]), .out(
        \mat_kron/mult_40_G2_G2_G1/B_not [7]) );
  inv \mat_kron/mult_40_G2_G2_G1/AN1_6_0  ( .in(\mat_add/r102/B_AS [6]), .out(
        \mat_kron/mult_40_G2_G2_G1/B_not [6]) );
  inv \mat_kron/mult_40_G2_G2_G1/AN1_5_0  ( .in(\mat_add/r102/B_AS [5]), .out(
        \mat_kron/mult_40_G2_G2_G1/B_not [5]) );
  inv \mat_kron/mult_40_G2_G2_G1/AN1_4_0  ( .in(\mat_add/r102/B_AS [4]), .out(
        \mat_kron/mult_40_G2_G2_G1/B_not [4]) );
  inv \mat_kron/mult_40_G2_G2_G1/AN1_3_0  ( .in(\mat_add/r102/B_AS [3]), .out(
        \mat_kron/mult_40_G2_G2_G1/B_not [3]) );
  inv \mat_kron/mult_40_G2_G2_G1/AN1_2_0  ( .in(\mat_add/r102/B_AS [2]), .out(
        \mat_kron/mult_40_G2_G2_G1/B_not [2]) );
  inv \mat_kron/mult_40_G2_G2_G1/AN1_1_0  ( .in(\mat_add/r102/B_AS [1]), .out(
        \mat_kron/mult_40_G2_G2_G1/B_not [1]) );
  inv \mat_kron/mult_40_G2_G2_G1/AN1_0_0  ( .in(\mat_add/r102/B_AS [0]), .out(
        \mat_kron/mult_40_G2_G2_G1/B_notx[0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN3_7_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [7]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[7][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_6_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [6]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[6][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_6_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [6]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[6][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_5_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[5][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_5_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[5][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_5_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[5][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_4_3  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[4][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_4_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[4][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_4_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[4][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_4_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[4][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_3_4  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[3][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_3_3  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[3][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_3_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[3][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_3_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[3][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_3_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[3][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_2_5  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[2][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_2_4  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[2][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_2_3  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[2][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_2_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[2][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_2_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[2][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_2_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[2][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_1_6  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [6]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[1][6] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_1_5  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[1][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_1_4  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[1][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_1_3  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[1][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_1_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[1][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_1_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[1][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_1_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[1][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN2_0_7  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [7]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[0][7] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_0_6  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [6]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[0][6] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_0_5  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[0][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_0_4  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[0][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_0_3  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[0][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_0_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[0][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_0_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1/ab[0][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1/AN1_0_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1/B_notx[0] ), .out(m_kro[72]) );
  inv \mat_kron/mult_40_G2_G2_G2_G1/AN1_7  ( .in(A[23]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [7]) );
  inv \mat_kron/mult_40_G2_G2_G2_G1/AN1_6  ( .in(A[22]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [6]) );
  inv \mat_kron/mult_40_G2_G2_G2_G1/AN1_5  ( .in(A[21]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [5]) );
  inv \mat_kron/mult_40_G2_G2_G2_G1/AN1_4  ( .in(A[20]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [4]) );
  inv \mat_kron/mult_40_G2_G2_G2_G1/AN1_3  ( .in(A[19]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [3]) );
  inv \mat_kron/mult_40_G2_G2_G2_G1/AN1_2  ( .in(A[18]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [2]) );
  inv \mat_kron/mult_40_G2_G2_G2_G1/AN1_1  ( .in(A[17]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [1]) );
  inv \mat_kron/mult_40_G2_G2_G2_G1/AN1_0  ( .in(A[16]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/A_notx[0] ) );
  inv \mat_kron/mult_40_G2_G2_G2_G1/AN1_7_0  ( .in(\mat_add/r106/B_AS [7]), 
        .out(\mat_kron/mult_40_G2_G2_G2_G1/B_not [7]) );
  inv \mat_kron/mult_40_G2_G2_G2_G1/AN1_6_0  ( .in(\mat_add/r106/B_AS [6]), 
        .out(\mat_kron/mult_40_G2_G2_G2_G1/B_not [6]) );
  inv \mat_kron/mult_40_G2_G2_G2_G1/AN1_5_0  ( .in(\mat_add/r106/B_AS [5]), 
        .out(\mat_kron/mult_40_G2_G2_G2_G1/B_not [5]) );
  inv \mat_kron/mult_40_G2_G2_G2_G1/AN1_4_0  ( .in(\mat_add/r106/B_AS [4]), 
        .out(\mat_kron/mult_40_G2_G2_G2_G1/B_not [4]) );
  inv \mat_kron/mult_40_G2_G2_G2_G1/AN1_3_0  ( .in(\mat_add/r106/B_AS [3]), 
        .out(\mat_kron/mult_40_G2_G2_G2_G1/B_not [3]) );
  inv \mat_kron/mult_40_G2_G2_G2_G1/AN1_2_0  ( .in(\mat_add/r106/B_AS [2]), 
        .out(\mat_kron/mult_40_G2_G2_G2_G1/B_not [2]) );
  inv \mat_kron/mult_40_G2_G2_G2_G1/AN1_1_0  ( .in(\mat_add/r106/B_AS [1]), 
        .out(\mat_kron/mult_40_G2_G2_G2_G1/B_not [1]) );
  inv \mat_kron/mult_40_G2_G2_G2_G1/AN1_0_0  ( .in(\mat_add/r106/B_AS [0]), 
        .out(\mat_kron/mult_40_G2_G2_G2_G1/B_notx[0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN3_7_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [7]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[7][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_6_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [6]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[6][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_6_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [6]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[6][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_5_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[5][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_5_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[5][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_5_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[5][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_4_3  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[4][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_4_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[4][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_4_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[4][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_4_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[4][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_3_4  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[3][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_3_3  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[3][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_3_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[3][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_3_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[3][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_3_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[3][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_2_5  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[2][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_2_4  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[2][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_2_3  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[2][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_2_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[2][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_2_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[2][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_2_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[2][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_1_6  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [6]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[1][6] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_1_5  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[1][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_1_4  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[1][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_1_3  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[1][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_1_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[1][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_1_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[1][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_1_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[1][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN2_0_7  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [7]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[0][7] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_0_6  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [6]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[0][6] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_0_5  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[0][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_0_4  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[0][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_0_3  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[0][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_0_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[0][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_0_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[0][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G1/AN1_0_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G1/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/B_notx[0] ), .out(m_kro[64]) );
  inv \mat_kron/mult_40_G2/AN1_7  ( .in(A[15]), .out(
        \mat_kron/mult_40_G2/A_not [7]) );
  inv \mat_kron/mult_40_G2/AN1_6  ( .in(A[14]), .out(
        \mat_kron/mult_40_G2/A_not [6]) );
  inv \mat_kron/mult_40_G2/AN1_5  ( .in(A[13]), .out(
        \mat_kron/mult_40_G2/A_not [5]) );
  inv \mat_kron/mult_40_G2/AN1_4  ( .in(A[12]), .out(
        \mat_kron/mult_40_G2/A_not [4]) );
  inv \mat_kron/mult_40_G2/AN1_3  ( .in(A[11]), .out(
        \mat_kron/mult_40_G2/A_not [3]) );
  inv \mat_kron/mult_40_G2/AN1_2  ( .in(A[10]), .out(
        \mat_kron/mult_40_G2/A_not [2]) );
  inv \mat_kron/mult_40_G2/AN1_1  ( .in(A[9]), .out(
        \mat_kron/mult_40_G2/A_not [1]) );
  inv \mat_kron/mult_40_G2/AN1_0  ( .in(A[8]), .out(
        \mat_kron/mult_40_G2/A_notx[0] ) );
  inv \mat_kron/mult_40_G2/AN1_7_0  ( .in(\mat_add/r94/B_AS [7]), .out(
        \mat_kron/mult_40_G2/B_not [7]) );
  inv \mat_kron/mult_40_G2/AN1_6_0  ( .in(\mat_add/r94/B_AS [6]), .out(
        \mat_kron/mult_40_G2/B_not [6]) );
  inv \mat_kron/mult_40_G2/AN1_5_0  ( .in(\mat_add/r94/B_AS [5]), .out(
        \mat_kron/mult_40_G2/B_not [5]) );
  inv \mat_kron/mult_40_G2/AN1_4_0  ( .in(\mat_add/r94/B_AS [4]), .out(
        \mat_kron/mult_40_G2/B_not [4]) );
  inv \mat_kron/mult_40_G2/AN1_3_0  ( .in(\mat_add/r94/B_AS [3]), .out(
        \mat_kron/mult_40_G2/B_not [3]) );
  inv \mat_kron/mult_40_G2/AN1_2_0  ( .in(\mat_add/r94/B_AS [2]), .out(
        \mat_kron/mult_40_G2/B_not [2]) );
  inv \mat_kron/mult_40_G2/AN1_1_0  ( .in(\mat_add/r94/B_AS [1]), .out(
        \mat_kron/mult_40_G2/B_not [1]) );
  inv \mat_kron/mult_40_G2/AN1_0_0  ( .in(\mat_add/r94/B_AS [0]), .out(
        \mat_kron/mult_40_G2/B_notx[0] ) );
  nor2 \mat_kron/mult_40_G2/AN3_7_0  ( .a(\mat_kron/mult_40_G2/A_not [7]), .b(
        \mat_kron/mult_40_G2/B_notx[0] ), .out(\mat_kron/mult_40_G2/ab[7][0] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_6_1  ( .a(\mat_kron/mult_40_G2/A_not [6]), .b(
        \mat_kron/mult_40_G2/B_not [1]), .out(\mat_kron/mult_40_G2/ab[6][1] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_6_0_0  ( .a(\mat_kron/mult_40_G2/A_not [6]), 
        .b(\mat_kron/mult_40_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2/ab[6][0] ) );
  nor2 \mat_kron/mult_40_G2/AN1_5_2  ( .a(\mat_kron/mult_40_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2/B_not [2]), .out(\mat_kron/mult_40_G2/ab[5][2] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_5_1  ( .a(\mat_kron/mult_40_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2/B_not [1]), .out(\mat_kron/mult_40_G2/ab[5][1] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_5_0_0  ( .a(\mat_kron/mult_40_G2/A_not [5]), 
        .b(\mat_kron/mult_40_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2/ab[5][0] ) );
  nor2 \mat_kron/mult_40_G2/AN1_4_3  ( .a(\mat_kron/mult_40_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2/B_not [3]), .out(\mat_kron/mult_40_G2/ab[4][3] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_4_2  ( .a(\mat_kron/mult_40_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2/B_not [2]), .out(\mat_kron/mult_40_G2/ab[4][2] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_4_1  ( .a(\mat_kron/mult_40_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2/B_not [1]), .out(\mat_kron/mult_40_G2/ab[4][1] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_4_0_0  ( .a(\mat_kron/mult_40_G2/A_not [4]), 
        .b(\mat_kron/mult_40_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2/ab[4][0] ) );
  nor2 \mat_kron/mult_40_G2/AN1_3_4  ( .a(\mat_kron/mult_40_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2/B_not [4]), .out(\mat_kron/mult_40_G2/ab[3][4] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_3_3  ( .a(\mat_kron/mult_40_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2/B_not [3]), .out(\mat_kron/mult_40_G2/ab[3][3] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_3_2  ( .a(\mat_kron/mult_40_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2/B_not [2]), .out(\mat_kron/mult_40_G2/ab[3][2] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_3_1  ( .a(\mat_kron/mult_40_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2/B_not [1]), .out(\mat_kron/mult_40_G2/ab[3][1] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_3_0_0  ( .a(\mat_kron/mult_40_G2/A_not [3]), 
        .b(\mat_kron/mult_40_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2/ab[3][0] ) );
  nor2 \mat_kron/mult_40_G2/AN1_2_5  ( .a(\mat_kron/mult_40_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2/B_not [5]), .out(\mat_kron/mult_40_G2/ab[2][5] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_2_4  ( .a(\mat_kron/mult_40_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2/B_not [4]), .out(\mat_kron/mult_40_G2/ab[2][4] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_2_3  ( .a(\mat_kron/mult_40_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2/B_not [3]), .out(\mat_kron/mult_40_G2/ab[2][3] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_2_2  ( .a(\mat_kron/mult_40_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2/B_not [2]), .out(\mat_kron/mult_40_G2/ab[2][2] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_2_1  ( .a(\mat_kron/mult_40_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2/B_not [1]), .out(\mat_kron/mult_40_G2/ab[2][1] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_2_0_0  ( .a(\mat_kron/mult_40_G2/A_not [2]), 
        .b(\mat_kron/mult_40_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2/ab[2][0] ) );
  nor2 \mat_kron/mult_40_G2/AN1_1_6  ( .a(\mat_kron/mult_40_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2/B_not [6]), .out(\mat_kron/mult_40_G2/ab[1][6] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_1_5  ( .a(\mat_kron/mult_40_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2/B_not [5]), .out(\mat_kron/mult_40_G2/ab[1][5] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_1_4  ( .a(\mat_kron/mult_40_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2/B_not [4]), .out(\mat_kron/mult_40_G2/ab[1][4] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_1_3  ( .a(\mat_kron/mult_40_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2/B_not [3]), .out(\mat_kron/mult_40_G2/ab[1][3] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_1_2  ( .a(\mat_kron/mult_40_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2/B_not [2]), .out(\mat_kron/mult_40_G2/ab[1][2] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_1_1  ( .a(\mat_kron/mult_40_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2/B_not [1]), .out(\mat_kron/mult_40_G2/ab[1][1] )
         );
  nor2 \mat_kron/mult_40_G2/AN1_1_0_0  ( .a(\mat_kron/mult_40_G2/A_not [1]), 
        .b(\mat_kron/mult_40_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2/ab[1][0] ) );
  nor2 \mat_kron/mult_40_G2/AN2_0_7  ( .a(\mat_kron/mult_40_G2/A_notx[0] ), 
        .b(\mat_kron/mult_40_G2/B_not [7]), .out(
        \mat_kron/mult_40_G2/ab[0][7] ) );
  nor2 \mat_kron/mult_40_G2/AN1_0_6  ( .a(\mat_kron/mult_40_G2/A_notx[0] ), 
        .b(\mat_kron/mult_40_G2/B_not [6]), .out(
        \mat_kron/mult_40_G2/ab[0][6] ) );
  nor2 \mat_kron/mult_40_G2/AN1_0_5  ( .a(\mat_kron/mult_40_G2/A_notx[0] ), 
        .b(\mat_kron/mult_40_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2/ab[0][5] ) );
  nor2 \mat_kron/mult_40_G2/AN1_0_4  ( .a(\mat_kron/mult_40_G2/A_notx[0] ), 
        .b(\mat_kron/mult_40_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2/ab[0][4] ) );
  nor2 \mat_kron/mult_40_G2/AN1_0_3  ( .a(\mat_kron/mult_40_G2/A_notx[0] ), 
        .b(\mat_kron/mult_40_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2/ab[0][3] ) );
  nor2 \mat_kron/mult_40_G2/AN1_0_2  ( .a(\mat_kron/mult_40_G2/A_notx[0] ), 
        .b(\mat_kron/mult_40_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2/ab[0][2] ) );
  nor2 \mat_kron/mult_40_G2/AN1_0_1  ( .a(\mat_kron/mult_40_G2/A_notx[0] ), 
        .b(\mat_kron/mult_40_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2/ab[0][1] ) );
  nor2 \mat_kron/mult_40_G2/AN1_0_0_0  ( .a(\mat_kron/mult_40_G2/A_notx[0] ), 
        .b(\mat_kron/mult_40_G2/B_notx[0] ), .out(m_kro[56]) );
  inv \mat_kron/mult_40_G2_G1_G1_G2/AN1_7  ( .in(A[15]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [7]) );
  inv \mat_kron/mult_40_G2_G1_G1_G2/AN1_6  ( .in(A[14]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [6]) );
  inv \mat_kron/mult_40_G2_G1_G1_G2/AN1_5  ( .in(A[13]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [5]) );
  inv \mat_kron/mult_40_G2_G1_G1_G2/AN1_4  ( .in(A[12]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [4]) );
  inv \mat_kron/mult_40_G2_G1_G1_G2/AN1_3  ( .in(A[11]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [3]) );
  inv \mat_kron/mult_40_G2_G1_G1_G2/AN1_2  ( .in(A[10]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [2]) );
  inv \mat_kron/mult_40_G2_G1_G1_G2/AN1_1  ( .in(A[9]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [1]) );
  inv \mat_kron/mult_40_G2_G1_G1_G2/AN1_0  ( .in(A[8]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/A_notx[0] ) );
  inv \mat_kron/mult_40_G2_G1_G1_G2/AN1_7_0  ( .in(\mat_add/r98/B_AS [7]), 
        .out(\mat_kron/mult_40_G2_G1_G1_G2/B_not [7]) );
  inv \mat_kron/mult_40_G2_G1_G1_G2/AN1_6_0  ( .in(\mat_add/r98/B_AS [6]), 
        .out(\mat_kron/mult_40_G2_G1_G1_G2/B_not [6]) );
  inv \mat_kron/mult_40_G2_G1_G1_G2/AN1_5_0  ( .in(\mat_add/r98/B_AS [5]), 
        .out(\mat_kron/mult_40_G2_G1_G1_G2/B_not [5]) );
  inv \mat_kron/mult_40_G2_G1_G1_G2/AN1_4_0  ( .in(\mat_add/r98/B_AS [4]), 
        .out(\mat_kron/mult_40_G2_G1_G1_G2/B_not [4]) );
  inv \mat_kron/mult_40_G2_G1_G1_G2/AN1_3_0  ( .in(\mat_add/r98/B_AS [3]), 
        .out(\mat_kron/mult_40_G2_G1_G1_G2/B_not [3]) );
  inv \mat_kron/mult_40_G2_G1_G1_G2/AN1_2_0  ( .in(\mat_add/r98/B_AS [2]), 
        .out(\mat_kron/mult_40_G2_G1_G1_G2/B_not [2]) );
  inv \mat_kron/mult_40_G2_G1_G1_G2/AN1_1_0  ( .in(\mat_add/r98/B_AS [1]), 
        .out(\mat_kron/mult_40_G2_G1_G1_G2/B_not [1]) );
  inv \mat_kron/mult_40_G2_G1_G1_G2/AN1_0_0  ( .in(\mat_add/r98/B_AS [0]), 
        .out(\mat_kron/mult_40_G2_G1_G1_G2/B_notx[0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN3_7_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [7]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[7][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_6_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [6]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[6][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_6_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [6]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[6][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_5_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[5][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_5_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[5][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_5_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[5][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_4_3  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[4][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_4_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[4][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_4_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[4][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_4_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[4][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_3_4  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[3][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_3_3  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[3][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_3_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[3][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_3_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[3][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_3_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[3][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_2_5  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[2][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_2_4  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[2][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_2_3  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[2][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_2_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[2][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_2_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[2][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_2_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[2][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_1_6  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [6]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[1][6] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_1_5  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[1][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_1_4  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[1][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_1_3  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[1][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_1_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[1][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_1_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[1][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_1_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[1][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN2_0_7  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [7]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[0][7] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_0_6  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [6]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[0][6] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_0_5  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[0][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_0_4  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[0][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_0_3  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[0][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_0_2  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[0][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_0_1  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[0][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G1_G2/AN1_0_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/B_notx[0] ), .out(m_kro[48]) );
  inv \mat_kron/mult_40_G2_G1_G2/AN1_7  ( .in(A[15]), .out(
        \mat_kron/mult_40_G2_G1_G2/A_not [7]) );
  inv \mat_kron/mult_40_G2_G1_G2/AN1_6  ( .in(A[14]), .out(
        \mat_kron/mult_40_G2_G1_G2/A_not [6]) );
  inv \mat_kron/mult_40_G2_G1_G2/AN1_5  ( .in(A[13]), .out(
        \mat_kron/mult_40_G2_G1_G2/A_not [5]) );
  inv \mat_kron/mult_40_G2_G1_G2/AN1_4  ( .in(A[12]), .out(
        \mat_kron/mult_40_G2_G1_G2/A_not [4]) );
  inv \mat_kron/mult_40_G2_G1_G2/AN1_3  ( .in(A[11]), .out(
        \mat_kron/mult_40_G2_G1_G2/A_not [3]) );
  inv \mat_kron/mult_40_G2_G1_G2/AN1_2  ( .in(A[10]), .out(
        \mat_kron/mult_40_G2_G1_G2/A_not [2]) );
  inv \mat_kron/mult_40_G2_G1_G2/AN1_1  ( .in(A[9]), .out(
        \mat_kron/mult_40_G2_G1_G2/A_not [1]) );
  inv \mat_kron/mult_40_G2_G1_G2/AN1_0  ( .in(A[8]), .out(
        \mat_kron/mult_40_G2_G1_G2/A_notx[0] ) );
  inv \mat_kron/mult_40_G2_G1_G2/AN1_7_0  ( .in(\mat_add/r102/B_AS [7]), .out(
        \mat_kron/mult_40_G2_G1_G2/B_not [7]) );
  inv \mat_kron/mult_40_G2_G1_G2/AN1_6_0  ( .in(\mat_add/r102/B_AS [6]), .out(
        \mat_kron/mult_40_G2_G1_G2/B_not [6]) );
  inv \mat_kron/mult_40_G2_G1_G2/AN1_5_0  ( .in(\mat_add/r102/B_AS [5]), .out(
        \mat_kron/mult_40_G2_G1_G2/B_not [5]) );
  inv \mat_kron/mult_40_G2_G1_G2/AN1_4_0  ( .in(\mat_add/r102/B_AS [4]), .out(
        \mat_kron/mult_40_G2_G1_G2/B_not [4]) );
  inv \mat_kron/mult_40_G2_G1_G2/AN1_3_0  ( .in(\mat_add/r102/B_AS [3]), .out(
        \mat_kron/mult_40_G2_G1_G2/B_not [3]) );
  inv \mat_kron/mult_40_G2_G1_G2/AN1_2_0  ( .in(\mat_add/r102/B_AS [2]), .out(
        \mat_kron/mult_40_G2_G1_G2/B_not [2]) );
  inv \mat_kron/mult_40_G2_G1_G2/AN1_1_0  ( .in(\mat_add/r102/B_AS [1]), .out(
        \mat_kron/mult_40_G2_G1_G2/B_not [1]) );
  inv \mat_kron/mult_40_G2_G1_G2/AN1_0_0  ( .in(\mat_add/r102/B_AS [0]), .out(
        \mat_kron/mult_40_G2_G1_G2/B_notx[0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN3_7_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [7]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[7][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_6_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [6]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[6][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_6_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [6]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[6][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_5_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[5][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_5_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[5][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_5_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[5][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_4_3  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[4][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_4_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[4][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_4_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[4][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_4_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[4][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_3_4  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[3][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_3_3  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[3][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_3_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[3][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_3_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[3][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_3_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[3][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_2_5  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[2][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_2_4  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[2][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_2_3  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[2][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_2_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[2][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_2_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[2][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_2_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[2][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_1_6  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [6]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[1][6] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_1_5  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[1][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_1_4  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[1][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_1_3  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[1][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_1_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[1][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_1_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[1][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_1_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[1][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN2_0_7  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [7]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[0][7] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_0_6  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [6]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[0][6] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_0_5  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[0][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_0_4  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[0][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_0_3  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[0][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_0_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[0][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_0_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2/ab[0][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2/AN1_0_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2/B_notx[0] ), .out(m_kro[24]) );
  inv \mat_kron/mult_40_G2_G2_G1_G2/AN1_7  ( .in(A[15]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [7]) );
  inv \mat_kron/mult_40_G2_G2_G1_G2/AN1_6  ( .in(A[14]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [6]) );
  inv \mat_kron/mult_40_G2_G2_G1_G2/AN1_5  ( .in(A[13]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [5]) );
  inv \mat_kron/mult_40_G2_G2_G1_G2/AN1_4  ( .in(A[12]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [4]) );
  inv \mat_kron/mult_40_G2_G2_G1_G2/AN1_3  ( .in(A[11]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [3]) );
  inv \mat_kron/mult_40_G2_G2_G1_G2/AN1_2  ( .in(A[10]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [2]) );
  inv \mat_kron/mult_40_G2_G2_G1_G2/AN1_1  ( .in(A[9]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [1]) );
  inv \mat_kron/mult_40_G2_G2_G1_G2/AN1_0  ( .in(A[8]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/A_notx[0] ) );
  inv \mat_kron/mult_40_G2_G2_G1_G2/AN1_7_0  ( .in(\mat_add/r106/B_AS [7]), 
        .out(\mat_kron/mult_40_G2_G2_G1_G2/B_not [7]) );
  inv \mat_kron/mult_40_G2_G2_G1_G2/AN1_6_0  ( .in(\mat_add/r106/B_AS [6]), 
        .out(\mat_kron/mult_40_G2_G2_G1_G2/B_not [6]) );
  inv \mat_kron/mult_40_G2_G2_G1_G2/AN1_5_0  ( .in(\mat_add/r106/B_AS [5]), 
        .out(\mat_kron/mult_40_G2_G2_G1_G2/B_not [5]) );
  inv \mat_kron/mult_40_G2_G2_G1_G2/AN1_4_0  ( .in(\mat_add/r106/B_AS [4]), 
        .out(\mat_kron/mult_40_G2_G2_G1_G2/B_not [4]) );
  inv \mat_kron/mult_40_G2_G2_G1_G2/AN1_3_0  ( .in(\mat_add/r106/B_AS [3]), 
        .out(\mat_kron/mult_40_G2_G2_G1_G2/B_not [3]) );
  inv \mat_kron/mult_40_G2_G2_G1_G2/AN1_2_0  ( .in(\mat_add/r106/B_AS [2]), 
        .out(\mat_kron/mult_40_G2_G2_G1_G2/B_not [2]) );
  inv \mat_kron/mult_40_G2_G2_G1_G2/AN1_1_0  ( .in(\mat_add/r106/B_AS [1]), 
        .out(\mat_kron/mult_40_G2_G2_G1_G2/B_not [1]) );
  inv \mat_kron/mult_40_G2_G2_G1_G2/AN1_0_0  ( .in(\mat_add/r106/B_AS [0]), 
        .out(\mat_kron/mult_40_G2_G2_G1_G2/B_notx[0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN3_7_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [7]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[7][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_6_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [6]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[6][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_6_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [6]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[6][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_5_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[5][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_5_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[5][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_5_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[5][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_4_3  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[4][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_4_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[4][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_4_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[4][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_4_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[4][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_3_4  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[3][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_3_3  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[3][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_3_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[3][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_3_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[3][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_3_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[3][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_2_5  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[2][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_2_4  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[2][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_2_3  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[2][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_2_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[2][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_2_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[2][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_2_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[2][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_1_6  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [6]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[1][6] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_1_5  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[1][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_1_4  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[1][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_1_3  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[1][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_1_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[1][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_1_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[1][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_1_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[1][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN2_0_7  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [7]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[0][7] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_0_6  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [6]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[0][6] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_0_5  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[0][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_0_4  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[0][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_0_3  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[0][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_0_2  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[0][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_0_1  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[0][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G1_G2/AN1_0_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G1_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/B_notx[0] ), .out(m_kro[16]) );
  inv \mat_kron/mult_40_G2_G2/AN1_7  ( .in(A[7]), .out(
        \mat_kron/mult_40_G2_G2/A_not [7]) );
  inv \mat_kron/mult_40_G2_G2/AN1_6  ( .in(A[6]), .out(
        \mat_kron/mult_40_G2_G2/A_not [6]) );
  inv \mat_kron/mult_40_G2_G2/AN1_5  ( .in(A[5]), .out(
        \mat_kron/mult_40_G2_G2/A_not [5]) );
  inv \mat_kron/mult_40_G2_G2/AN1_4  ( .in(A[4]), .out(
        \mat_kron/mult_40_G2_G2/A_not [4]) );
  inv \mat_kron/mult_40_G2_G2/AN1_3  ( .in(A[3]), .out(
        \mat_kron/mult_40_G2_G2/A_not [3]) );
  inv \mat_kron/mult_40_G2_G2/AN1_2  ( .in(A[2]), .out(
        \mat_kron/mult_40_G2_G2/A_not [2]) );
  inv \mat_kron/mult_40_G2_G2/AN1_1  ( .in(A[1]), .out(
        \mat_kron/mult_40_G2_G2/A_not [1]) );
  inv \mat_kron/mult_40_G2_G2/AN1_0  ( .in(A[0]), .out(
        \mat_kron/mult_40_G2_G2/A_notx[0] ) );
  inv \mat_kron/mult_40_G2_G2/AN1_7_0  ( .in(\mat_add/r94/B_AS [7]), .out(
        \mat_kron/mult_40_G2_G2/B_not [7]) );
  inv \mat_kron/mult_40_G2_G2/AN1_6_0  ( .in(\mat_add/r94/B_AS [6]), .out(
        \mat_kron/mult_40_G2_G2/B_not [6]) );
  inv \mat_kron/mult_40_G2_G2/AN1_5_0  ( .in(\mat_add/r94/B_AS [5]), .out(
        \mat_kron/mult_40_G2_G2/B_not [5]) );
  inv \mat_kron/mult_40_G2_G2/AN1_4_0  ( .in(\mat_add/r94/B_AS [4]), .out(
        \mat_kron/mult_40_G2_G2/B_not [4]) );
  inv \mat_kron/mult_40_G2_G2/AN1_3_0  ( .in(\mat_add/r94/B_AS [3]), .out(
        \mat_kron/mult_40_G2_G2/B_not [3]) );
  inv \mat_kron/mult_40_G2_G2/AN1_2_0  ( .in(\mat_add/r94/B_AS [2]), .out(
        \mat_kron/mult_40_G2_G2/B_not [2]) );
  inv \mat_kron/mult_40_G2_G2/AN1_1_0  ( .in(\mat_add/r94/B_AS [1]), .out(
        \mat_kron/mult_40_G2_G2/B_not [1]) );
  inv \mat_kron/mult_40_G2_G2/AN1_0_0  ( .in(\mat_add/r94/B_AS [0]), .out(
        \mat_kron/mult_40_G2_G2/B_notx[0] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN3_7_0  ( .a(\mat_kron/mult_40_G2_G2/A_not [7]), .b(\mat_kron/mult_40_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2/ab[7][0] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_6_1  ( .a(\mat_kron/mult_40_G2_G2/A_not [6]), .b(\mat_kron/mult_40_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2/ab[6][1] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_6_0_0  ( .a(
        \mat_kron/mult_40_G2_G2/A_not [6]), .b(
        \mat_kron/mult_40_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2/ab[6][0] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_5_2  ( .a(\mat_kron/mult_40_G2_G2/A_not [5]), .b(\mat_kron/mult_40_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2/ab[5][2] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_5_1  ( .a(\mat_kron/mult_40_G2_G2/A_not [5]), .b(\mat_kron/mult_40_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2/ab[5][1] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_5_0_0  ( .a(
        \mat_kron/mult_40_G2_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2/ab[5][0] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_4_3  ( .a(\mat_kron/mult_40_G2_G2/A_not [4]), .b(\mat_kron/mult_40_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2/ab[4][3] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_4_2  ( .a(\mat_kron/mult_40_G2_G2/A_not [4]), .b(\mat_kron/mult_40_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2/ab[4][2] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_4_1  ( .a(\mat_kron/mult_40_G2_G2/A_not [4]), .b(\mat_kron/mult_40_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2/ab[4][1] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_4_0_0  ( .a(
        \mat_kron/mult_40_G2_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2/ab[4][0] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_3_4  ( .a(\mat_kron/mult_40_G2_G2/A_not [3]), .b(\mat_kron/mult_40_G2_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2/ab[3][4] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_3_3  ( .a(\mat_kron/mult_40_G2_G2/A_not [3]), .b(\mat_kron/mult_40_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2/ab[3][3] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_3_2  ( .a(\mat_kron/mult_40_G2_G2/A_not [3]), .b(\mat_kron/mult_40_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2/ab[3][2] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_3_1  ( .a(\mat_kron/mult_40_G2_G2/A_not [3]), .b(\mat_kron/mult_40_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2/ab[3][1] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_3_0_0  ( .a(
        \mat_kron/mult_40_G2_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2/ab[3][0] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_2_5  ( .a(\mat_kron/mult_40_G2_G2/A_not [2]), .b(\mat_kron/mult_40_G2_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2/ab[2][5] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_2_4  ( .a(\mat_kron/mult_40_G2_G2/A_not [2]), .b(\mat_kron/mult_40_G2_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2/ab[2][4] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_2_3  ( .a(\mat_kron/mult_40_G2_G2/A_not [2]), .b(\mat_kron/mult_40_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2/ab[2][3] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_2_2  ( .a(\mat_kron/mult_40_G2_G2/A_not [2]), .b(\mat_kron/mult_40_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2/ab[2][2] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_2_1  ( .a(\mat_kron/mult_40_G2_G2/A_not [2]), .b(\mat_kron/mult_40_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2/ab[2][1] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_2_0_0  ( .a(
        \mat_kron/mult_40_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2/ab[2][0] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_1_6  ( .a(\mat_kron/mult_40_G2_G2/A_not [1]), .b(\mat_kron/mult_40_G2_G2/B_not [6]), .out(
        \mat_kron/mult_40_G2_G2/ab[1][6] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_1_5  ( .a(\mat_kron/mult_40_G2_G2/A_not [1]), .b(\mat_kron/mult_40_G2_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2/ab[1][5] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_1_4  ( .a(\mat_kron/mult_40_G2_G2/A_not [1]), .b(\mat_kron/mult_40_G2_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2/ab[1][4] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_1_3  ( .a(\mat_kron/mult_40_G2_G2/A_not [1]), .b(\mat_kron/mult_40_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2/ab[1][3] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_1_2  ( .a(\mat_kron/mult_40_G2_G2/A_not [1]), .b(\mat_kron/mult_40_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2/ab[1][2] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_1_1  ( .a(\mat_kron/mult_40_G2_G2/A_not [1]), .b(\mat_kron/mult_40_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2/ab[1][1] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_1_0_0  ( .a(
        \mat_kron/mult_40_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2/ab[1][0] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN2_0_7  ( .a(
        \mat_kron/mult_40_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2/B_not [7]), .out(
        \mat_kron/mult_40_G2_G2/ab[0][7] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_0_6  ( .a(
        \mat_kron/mult_40_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2/B_not [6]), .out(
        \mat_kron/mult_40_G2_G2/ab[0][6] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_0_5  ( .a(
        \mat_kron/mult_40_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2/ab[0][5] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_0_4  ( .a(
        \mat_kron/mult_40_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2/ab[0][4] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_0_3  ( .a(
        \mat_kron/mult_40_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2/ab[0][3] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_0_2  ( .a(
        \mat_kron/mult_40_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2/ab[0][2] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_0_1  ( .a(
        \mat_kron/mult_40_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2/ab[0][1] ) );
  nor2 \mat_kron/mult_40_G2_G2/AN1_0_0_0  ( .a(
        \mat_kron/mult_40_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2/B_notx[0] ), .out(m_kro[40]) );
  inv \mat_kron/mult_40_G2_G1_G2_G2/AN1_7  ( .in(A[7]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [7]) );
  inv \mat_kron/mult_40_G2_G1_G2_G2/AN1_6  ( .in(A[6]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [6]) );
  inv \mat_kron/mult_40_G2_G1_G2_G2/AN1_5  ( .in(A[5]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [5]) );
  inv \mat_kron/mult_40_G2_G1_G2_G2/AN1_4  ( .in(A[4]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [4]) );
  inv \mat_kron/mult_40_G2_G1_G2_G2/AN1_3  ( .in(A[3]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [3]) );
  inv \mat_kron/mult_40_G2_G1_G2_G2/AN1_2  ( .in(A[2]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [2]) );
  inv \mat_kron/mult_40_G2_G1_G2_G2/AN1_1  ( .in(A[1]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [1]) );
  inv \mat_kron/mult_40_G2_G1_G2_G2/AN1_0  ( .in(A[0]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/A_notx[0] ) );
  inv \mat_kron/mult_40_G2_G1_G2_G2/AN1_7_0  ( .in(\mat_add/r98/B_AS [7]), 
        .out(\mat_kron/mult_40_G2_G1_G2_G2/B_not [7]) );
  inv \mat_kron/mult_40_G2_G1_G2_G2/AN1_6_0  ( .in(\mat_add/r98/B_AS [6]), 
        .out(\mat_kron/mult_40_G2_G1_G2_G2/B_not [6]) );
  inv \mat_kron/mult_40_G2_G1_G2_G2/AN1_5_0  ( .in(\mat_add/r98/B_AS [5]), 
        .out(\mat_kron/mult_40_G2_G1_G2_G2/B_not [5]) );
  inv \mat_kron/mult_40_G2_G1_G2_G2/AN1_4_0  ( .in(\mat_add/r98/B_AS [4]), 
        .out(\mat_kron/mult_40_G2_G1_G2_G2/B_not [4]) );
  inv \mat_kron/mult_40_G2_G1_G2_G2/AN1_3_0  ( .in(\mat_add/r98/B_AS [3]), 
        .out(\mat_kron/mult_40_G2_G1_G2_G2/B_not [3]) );
  inv \mat_kron/mult_40_G2_G1_G2_G2/AN1_2_0  ( .in(\mat_add/r98/B_AS [2]), 
        .out(\mat_kron/mult_40_G2_G1_G2_G2/B_not [2]) );
  inv \mat_kron/mult_40_G2_G1_G2_G2/AN1_1_0  ( .in(\mat_add/r98/B_AS [1]), 
        .out(\mat_kron/mult_40_G2_G1_G2_G2/B_not [1]) );
  inv \mat_kron/mult_40_G2_G1_G2_G2/AN1_0_0  ( .in(\mat_add/r98/B_AS [0]), 
        .out(\mat_kron/mult_40_G2_G1_G2_G2/B_notx[0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN3_7_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [7]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[7][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_6_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [6]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[6][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_6_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [6]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[6][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_5_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[5][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_5_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[5][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_5_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[5][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_4_3  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[4][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_4_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[4][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_4_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[4][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_4_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[4][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_3_4  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[3][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_3_3  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[3][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_3_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[3][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_3_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[3][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_3_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[3][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_2_5  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[2][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_2_4  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[2][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_2_3  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[2][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_2_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[2][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_2_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[2][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_2_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[2][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_1_6  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [6]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[1][6] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_1_5  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[1][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_1_4  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[1][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_1_3  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[1][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_1_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[1][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_1_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[1][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_1_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[1][0] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN2_0_7  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [7]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[0][7] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_0_6  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [6]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[0][6] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_0_5  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[0][5] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_0_4  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[0][4] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_0_3  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[0][3] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_0_2  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[0][2] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_0_1  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[0][1] ) );
  nor2 \mat_kron/mult_40_G2_G1_G2_G2/AN1_0_0_0  ( .a(
        \mat_kron/mult_40_G2_G1_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/B_notx[0] ), .out(m_kro[32]) );
  inv \mat_kron/mult_40_G2_G2_G2/AN1_7  ( .in(A[7]), .out(
        \mat_kron/mult_40_G2_G2_G2/A_not [7]) );
  inv \mat_kron/mult_40_G2_G2_G2/AN1_6  ( .in(A[6]), .out(
        \mat_kron/mult_40_G2_G2_G2/A_not [6]) );
  inv \mat_kron/mult_40_G2_G2_G2/AN1_5  ( .in(A[5]), .out(
        \mat_kron/mult_40_G2_G2_G2/A_not [5]) );
  inv \mat_kron/mult_40_G2_G2_G2/AN1_4  ( .in(A[4]), .out(
        \mat_kron/mult_40_G2_G2_G2/A_not [4]) );
  inv \mat_kron/mult_40_G2_G2_G2/AN1_3  ( .in(A[3]), .out(
        \mat_kron/mult_40_G2_G2_G2/A_not [3]) );
  inv \mat_kron/mult_40_G2_G2_G2/AN1_2  ( .in(A[2]), .out(
        \mat_kron/mult_40_G2_G2_G2/A_not [2]) );
  inv \mat_kron/mult_40_G2_G2_G2/AN1_1  ( .in(A[1]), .out(
        \mat_kron/mult_40_G2_G2_G2/A_not [1]) );
  inv \mat_kron/mult_40_G2_G2_G2/AN1_0  ( .in(A[0]), .out(
        \mat_kron/mult_40_G2_G2_G2/A_notx[0] ) );
  inv \mat_kron/mult_40_G2_G2_G2/AN1_7_0  ( .in(\mat_add/r102/B_AS [7]), .out(
        \mat_kron/mult_40_G2_G2_G2/B_not [7]) );
  inv \mat_kron/mult_40_G2_G2_G2/AN1_6_0  ( .in(\mat_add/r102/B_AS [6]), .out(
        \mat_kron/mult_40_G2_G2_G2/B_not [6]) );
  inv \mat_kron/mult_40_G2_G2_G2/AN1_5_0  ( .in(\mat_add/r102/B_AS [5]), .out(
        \mat_kron/mult_40_G2_G2_G2/B_not [5]) );
  inv \mat_kron/mult_40_G2_G2_G2/AN1_4_0  ( .in(\mat_add/r102/B_AS [4]), .out(
        \mat_kron/mult_40_G2_G2_G2/B_not [4]) );
  inv \mat_kron/mult_40_G2_G2_G2/AN1_3_0  ( .in(\mat_add/r102/B_AS [3]), .out(
        \mat_kron/mult_40_G2_G2_G2/B_not [3]) );
  inv \mat_kron/mult_40_G2_G2_G2/AN1_2_0  ( .in(\mat_add/r102/B_AS [2]), .out(
        \mat_kron/mult_40_G2_G2_G2/B_not [2]) );
  inv \mat_kron/mult_40_G2_G2_G2/AN1_1_0  ( .in(\mat_add/r102/B_AS [1]), .out(
        \mat_kron/mult_40_G2_G2_G2/B_not [1]) );
  inv \mat_kron/mult_40_G2_G2_G2/AN1_0_0  ( .in(\mat_add/r102/B_AS [0]), .out(
        \mat_kron/mult_40_G2_G2_G2/B_notx[0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN3_7_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [7]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[7][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_6_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [6]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[6][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_6_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [6]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[6][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_5_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[5][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_5_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[5][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_5_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[5][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_4_3  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[4][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_4_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[4][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_4_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[4][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_4_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[4][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_3_4  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[3][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_3_3  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[3][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_3_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[3][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_3_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[3][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_3_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[3][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_2_5  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[2][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_2_4  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[2][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_2_3  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[2][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_2_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[2][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_2_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[2][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_2_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[2][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_1_6  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [6]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[1][6] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_1_5  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[1][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_1_4  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[1][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_1_3  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[1][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_1_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[1][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_1_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[1][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_1_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[1][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN2_0_7  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [7]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[0][7] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_0_6  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [6]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[0][6] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_0_5  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[0][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_0_4  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[0][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_0_3  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[0][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_0_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[0][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_0_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2/ab[0][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2/AN1_0_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2/B_notx[0] ), .out(m_kro[8]) );
  inv \mat_kron/mult_40_G2_G2_G2_G2/AN1_7  ( .in(A[7]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [7]) );
  inv \mat_kron/mult_40_G2_G2_G2_G2/AN1_6  ( .in(A[6]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [6]) );
  inv \mat_kron/mult_40_G2_G2_G2_G2/AN1_5  ( .in(A[5]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [5]) );
  inv \mat_kron/mult_40_G2_G2_G2_G2/AN1_4  ( .in(A[4]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [4]) );
  inv \mat_kron/mult_40_G2_G2_G2_G2/AN1_3  ( .in(A[3]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [3]) );
  inv \mat_kron/mult_40_G2_G2_G2_G2/AN1_2  ( .in(A[2]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [2]) );
  inv \mat_kron/mult_40_G2_G2_G2_G2/AN1_1  ( .in(A[1]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [1]) );
  inv \mat_kron/mult_40_G2_G2_G2_G2/AN1_0  ( .in(A[0]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/A_notx[0] ) );
  inv \mat_kron/mult_40_G2_G2_G2_G2/AN1_7_0  ( .in(\mat_add/r106/B_AS [7]), 
        .out(\mat_kron/mult_40_G2_G2_G2_G2/B_not [7]) );
  inv \mat_kron/mult_40_G2_G2_G2_G2/AN1_6_0  ( .in(\mat_add/r106/B_AS [6]), 
        .out(\mat_kron/mult_40_G2_G2_G2_G2/B_not [6]) );
  inv \mat_kron/mult_40_G2_G2_G2_G2/AN1_5_0  ( .in(\mat_add/r106/B_AS [5]), 
        .out(\mat_kron/mult_40_G2_G2_G2_G2/B_not [5]) );
  inv \mat_kron/mult_40_G2_G2_G2_G2/AN1_4_0  ( .in(\mat_add/r106/B_AS [4]), 
        .out(\mat_kron/mult_40_G2_G2_G2_G2/B_not [4]) );
  inv \mat_kron/mult_40_G2_G2_G2_G2/AN1_3_0  ( .in(\mat_add/r106/B_AS [3]), 
        .out(\mat_kron/mult_40_G2_G2_G2_G2/B_not [3]) );
  inv \mat_kron/mult_40_G2_G2_G2_G2/AN1_2_0  ( .in(\mat_add/r106/B_AS [2]), 
        .out(\mat_kron/mult_40_G2_G2_G2_G2/B_not [2]) );
  inv \mat_kron/mult_40_G2_G2_G2_G2/AN1_1_0  ( .in(\mat_add/r106/B_AS [1]), 
        .out(\mat_kron/mult_40_G2_G2_G2_G2/B_not [1]) );
  inv \mat_kron/mult_40_G2_G2_G2_G2/AN1_0_0  ( .in(\mat_add/r106/B_AS [0]), 
        .out(\mat_kron/mult_40_G2_G2_G2_G2/B_notx[0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN3_7_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [7]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[7][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_6_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [6]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[6][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_6_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [6]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[6][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_5_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[5][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_5_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[5][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_5_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [5]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[5][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_4_3  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[4][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_4_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[4][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_4_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[4][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_4_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [4]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[4][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_3_4  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[3][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_3_3  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[3][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_3_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[3][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_3_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[3][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_3_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [3]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[3][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_2_5  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[2][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_2_4  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[2][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_2_3  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[2][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_2_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[2][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_2_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[2][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_2_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [2]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[2][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_1_6  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [6]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[1][6] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_1_5  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[1][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_1_4  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[1][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_1_3  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[1][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_1_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[1][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_1_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[1][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_1_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_not [1]), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_notx[0] ), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[1][0] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN2_0_7  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [7]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[0][7] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_0_6  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [6]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[0][6] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_0_5  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [5]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[0][5] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_0_4  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [4]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[0][4] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_0_3  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [3]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[0][3] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_0_2  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [2]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[0][2] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_0_1  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_not [1]), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[0][1] ) );
  nor2 \mat_kron/mult_40_G2_G2_G2_G2/AN1_0_0_0  ( .a(
        \mat_kron/mult_40_G2_G2_G2_G2/A_notx[0] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/B_notx[0] ), .out(m_kro[0]) );
  inv \mat_mul/mult_37/AN1_7  ( .in(A[31]), .out(\mat_mul/mult_37/A_not [7])
         );
  inv \mat_mul/mult_37/AN1_6  ( .in(A[30]), .out(\mat_mul/mult_37/A_not [6])
         );
  inv \mat_mul/mult_37/AN1_5  ( .in(A[29]), .out(\mat_mul/mult_37/A_not [5])
         );
  inv \mat_mul/mult_37/AN1_4  ( .in(A[28]), .out(\mat_mul/mult_37/A_not [4])
         );
  inv \mat_mul/mult_37/AN1_3  ( .in(A[27]), .out(\mat_mul/mult_37/A_not [3])
         );
  inv \mat_mul/mult_37/AN1_2  ( .in(A[26]), .out(\mat_mul/mult_37/A_not [2])
         );
  inv \mat_mul/mult_37/AN1_1  ( .in(A[25]), .out(\mat_mul/mult_37/A_not [1])
         );
  inv \mat_mul/mult_37/AN1_0  ( .in(A[24]), .out(\mat_mul/mult_37/A_notx[0] )
         );
  inv \mat_mul/mult_37/AN1_7_0  ( .in(\mat_add/r94/B_AS [7]), .out(
        \mat_mul/mult_37/B_not [7]) );
  inv \mat_mul/mult_37/AN1_6_0  ( .in(\mat_add/r94/B_AS [6]), .out(
        \mat_mul/mult_37/B_not [6]) );
  inv \mat_mul/mult_37/AN1_5_0  ( .in(\mat_add/r94/B_AS [5]), .out(
        \mat_mul/mult_37/B_not [5]) );
  inv \mat_mul/mult_37/AN1_4_0  ( .in(\mat_add/r94/B_AS [4]), .out(
        \mat_mul/mult_37/B_not [4]) );
  inv \mat_mul/mult_37/AN1_3_0  ( .in(\mat_add/r94/B_AS [3]), .out(
        \mat_mul/mult_37/B_not [3]) );
  inv \mat_mul/mult_37/AN1_2_0  ( .in(\mat_add/r94/B_AS [2]), .out(
        \mat_mul/mult_37/B_not [2]) );
  inv \mat_mul/mult_37/AN1_1_0  ( .in(\mat_add/r94/B_AS [1]), .out(
        \mat_mul/mult_37/B_not [1]) );
  inv \mat_mul/mult_37/AN1_0_0  ( .in(\mat_add/r94/B_AS [0]), .out(
        \mat_mul/mult_37/B_notx[0] ) );
  nor2 \mat_mul/mult_37/AN3_7_0  ( .a(\mat_mul/mult_37/A_not [7]), .b(
        \mat_mul/mult_37/B_notx[0] ), .out(\mat_mul/mult_37/ab[7][0] ) );
  nor2 \mat_mul/mult_37/AN1_6_1  ( .a(\mat_mul/mult_37/A_not [6]), .b(
        \mat_mul/mult_37/B_not [1]), .out(\mat_mul/mult_37/ab[6][1] ) );
  nor2 \mat_mul/mult_37/AN1_6_0_0  ( .a(\mat_mul/mult_37/A_not [6]), .b(
        \mat_mul/mult_37/B_notx[0] ), .out(\mat_mul/mult_37/ab[6][0] ) );
  nor2 \mat_mul/mult_37/AN1_5_2  ( .a(\mat_mul/mult_37/A_not [5]), .b(
        \mat_mul/mult_37/B_not [2]), .out(\mat_mul/mult_37/ab[5][2] ) );
  nor2 \mat_mul/mult_37/AN1_5_1  ( .a(\mat_mul/mult_37/A_not [5]), .b(
        \mat_mul/mult_37/B_not [1]), .out(\mat_mul/mult_37/ab[5][1] ) );
  nor2 \mat_mul/mult_37/AN1_5_0_0  ( .a(\mat_mul/mult_37/A_not [5]), .b(
        \mat_mul/mult_37/B_notx[0] ), .out(\mat_mul/mult_37/ab[5][0] ) );
  nor2 \mat_mul/mult_37/AN1_4_3  ( .a(\mat_mul/mult_37/A_not [4]), .b(
        \mat_mul/mult_37/B_not [3]), .out(\mat_mul/mult_37/ab[4][3] ) );
  nor2 \mat_mul/mult_37/AN1_4_2  ( .a(\mat_mul/mult_37/A_not [4]), .b(
        \mat_mul/mult_37/B_not [2]), .out(\mat_mul/mult_37/ab[4][2] ) );
  nor2 \mat_mul/mult_37/AN1_4_1  ( .a(\mat_mul/mult_37/A_not [4]), .b(
        \mat_mul/mult_37/B_not [1]), .out(\mat_mul/mult_37/ab[4][1] ) );
  nor2 \mat_mul/mult_37/AN1_4_0_0  ( .a(\mat_mul/mult_37/A_not [4]), .b(
        \mat_mul/mult_37/B_notx[0] ), .out(\mat_mul/mult_37/ab[4][0] ) );
  nor2 \mat_mul/mult_37/AN1_3_4  ( .a(\mat_mul/mult_37/A_not [3]), .b(
        \mat_mul/mult_37/B_not [4]), .out(\mat_mul/mult_37/ab[3][4] ) );
  nor2 \mat_mul/mult_37/AN1_3_3  ( .a(\mat_mul/mult_37/A_not [3]), .b(
        \mat_mul/mult_37/B_not [3]), .out(\mat_mul/mult_37/ab[3][3] ) );
  nor2 \mat_mul/mult_37/AN1_3_2  ( .a(\mat_mul/mult_37/A_not [3]), .b(
        \mat_mul/mult_37/B_not [2]), .out(\mat_mul/mult_37/ab[3][2] ) );
  nor2 \mat_mul/mult_37/AN1_3_1  ( .a(\mat_mul/mult_37/A_not [3]), .b(
        \mat_mul/mult_37/B_not [1]), .out(\mat_mul/mult_37/ab[3][1] ) );
  nor2 \mat_mul/mult_37/AN1_3_0_0  ( .a(\mat_mul/mult_37/A_not [3]), .b(
        \mat_mul/mult_37/B_notx[0] ), .out(\mat_mul/mult_37/ab[3][0] ) );
  nor2 \mat_mul/mult_37/AN1_2_5  ( .a(\mat_mul/mult_37/A_not [2]), .b(
        \mat_mul/mult_37/B_not [5]), .out(\mat_mul/mult_37/ab[2][5] ) );
  nor2 \mat_mul/mult_37/AN1_2_4  ( .a(\mat_mul/mult_37/A_not [2]), .b(
        \mat_mul/mult_37/B_not [4]), .out(\mat_mul/mult_37/ab[2][4] ) );
  nor2 \mat_mul/mult_37/AN1_2_3  ( .a(\mat_mul/mult_37/A_not [2]), .b(
        \mat_mul/mult_37/B_not [3]), .out(\mat_mul/mult_37/ab[2][3] ) );
  nor2 \mat_mul/mult_37/AN1_2_2  ( .a(\mat_mul/mult_37/A_not [2]), .b(
        \mat_mul/mult_37/B_not [2]), .out(\mat_mul/mult_37/ab[2][2] ) );
  nor2 \mat_mul/mult_37/AN1_2_1  ( .a(\mat_mul/mult_37/A_not [2]), .b(
        \mat_mul/mult_37/B_not [1]), .out(\mat_mul/mult_37/ab[2][1] ) );
  nor2 \mat_mul/mult_37/AN1_2_0_0  ( .a(\mat_mul/mult_37/A_not [2]), .b(
        \mat_mul/mult_37/B_notx[0] ), .out(\mat_mul/mult_37/ab[2][0] ) );
  nor2 \mat_mul/mult_37/AN1_1_6  ( .a(\mat_mul/mult_37/A_not [1]), .b(
        \mat_mul/mult_37/B_not [6]), .out(\mat_mul/mult_37/ab[1][6] ) );
  nor2 \mat_mul/mult_37/AN1_1_5  ( .a(\mat_mul/mult_37/A_not [1]), .b(
        \mat_mul/mult_37/B_not [5]), .out(\mat_mul/mult_37/ab[1][5] ) );
  nor2 \mat_mul/mult_37/AN1_1_4  ( .a(\mat_mul/mult_37/A_not [1]), .b(
        \mat_mul/mult_37/B_not [4]), .out(\mat_mul/mult_37/ab[1][4] ) );
  nor2 \mat_mul/mult_37/AN1_1_3  ( .a(\mat_mul/mult_37/A_not [1]), .b(
        \mat_mul/mult_37/B_not [3]), .out(\mat_mul/mult_37/ab[1][3] ) );
  nor2 \mat_mul/mult_37/AN1_1_2  ( .a(\mat_mul/mult_37/A_not [1]), .b(
        \mat_mul/mult_37/B_not [2]), .out(\mat_mul/mult_37/ab[1][2] ) );
  nor2 \mat_mul/mult_37/AN1_1_1  ( .a(\mat_mul/mult_37/A_not [1]), .b(
        \mat_mul/mult_37/B_not [1]), .out(\mat_mul/mult_37/ab[1][1] ) );
  nor2 \mat_mul/mult_37/AN1_1_0_0  ( .a(\mat_mul/mult_37/A_not [1]), .b(
        \mat_mul/mult_37/B_notx[0] ), .out(\mat_mul/mult_37/ab[1][0] ) );
  nor2 \mat_mul/mult_37/AN2_0_7  ( .a(\mat_mul/mult_37/A_notx[0] ), .b(
        \mat_mul/mult_37/B_not [7]), .out(\mat_mul/mult_37/ab[0][7] ) );
  nor2 \mat_mul/mult_37/AN1_0_6  ( .a(\mat_mul/mult_37/A_notx[0] ), .b(
        \mat_mul/mult_37/B_not [6]), .out(\mat_mul/mult_37/ab[0][6] ) );
  nor2 \mat_mul/mult_37/AN1_0_5  ( .a(\mat_mul/mult_37/A_notx[0] ), .b(
        \mat_mul/mult_37/B_not [5]), .out(\mat_mul/mult_37/ab[0][5] ) );
  nor2 \mat_mul/mult_37/AN1_0_4  ( .a(\mat_mul/mult_37/A_notx[0] ), .b(
        \mat_mul/mult_37/B_not [4]), .out(\mat_mul/mult_37/ab[0][4] ) );
  nor2 \mat_mul/mult_37/AN1_0_3  ( .a(\mat_mul/mult_37/A_notx[0] ), .b(
        \mat_mul/mult_37/B_not [3]), .out(\mat_mul/mult_37/ab[0][3] ) );
  nor2 \mat_mul/mult_37/AN1_0_2  ( .a(\mat_mul/mult_37/A_notx[0] ), .b(
        \mat_mul/mult_37/B_not [2]), .out(\mat_mul/mult_37/ab[0][2] ) );
  nor2 \mat_mul/mult_37/AN1_0_1  ( .a(\mat_mul/mult_37/A_notx[0] ), .b(
        \mat_mul/mult_37/B_not [1]), .out(\mat_mul/mult_37/ab[0][1] ) );
  nor2 \mat_mul/mult_37/AN1_0_0_0  ( .a(\mat_mul/mult_37/A_notx[0] ), .b(
        \mat_mul/mult_37/B_notx[0] ), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[0] ) );
  inv \mat_mul/mult_37_G2_G1_G1/AN1_7  ( .in(A[23]), .out(
        \mat_mul/mult_37_G2_G1_G1/A_not [7]) );
  inv \mat_mul/mult_37_G2_G1_G1/AN1_6  ( .in(A[22]), .out(
        \mat_mul/mult_37_G2_G1_G1/A_not [6]) );
  inv \mat_mul/mult_37_G2_G1_G1/AN1_5  ( .in(A[21]), .out(
        \mat_mul/mult_37_G2_G1_G1/A_not [5]) );
  inv \mat_mul/mult_37_G2_G1_G1/AN1_4  ( .in(A[20]), .out(
        \mat_mul/mult_37_G2_G1_G1/A_not [4]) );
  inv \mat_mul/mult_37_G2_G1_G1/AN1_3  ( .in(A[19]), .out(
        \mat_mul/mult_37_G2_G1_G1/A_not [3]) );
  inv \mat_mul/mult_37_G2_G1_G1/AN1_2  ( .in(A[18]), .out(
        \mat_mul/mult_37_G2_G1_G1/A_not [2]) );
  inv \mat_mul/mult_37_G2_G1_G1/AN1_1  ( .in(A[17]), .out(
        \mat_mul/mult_37_G2_G1_G1/A_not [1]) );
  inv \mat_mul/mult_37_G2_G1_G1/AN1_0  ( .in(A[16]), .out(
        \mat_mul/mult_37_G2_G1_G1/A_notx[0] ) );
  inv \mat_mul/mult_37_G2_G1_G1/AN1_7_0  ( .in(\mat_add/r102/B_AS [7]), .out(
        \mat_mul/mult_37_G2_G1_G1/B_not [7]) );
  inv \mat_mul/mult_37_G2_G1_G1/AN1_6_0  ( .in(\mat_add/r102/B_AS [6]), .out(
        \mat_mul/mult_37_G2_G1_G1/B_not [6]) );
  inv \mat_mul/mult_37_G2_G1_G1/AN1_5_0  ( .in(\mat_add/r102/B_AS [5]), .out(
        \mat_mul/mult_37_G2_G1_G1/B_not [5]) );
  inv \mat_mul/mult_37_G2_G1_G1/AN1_4_0  ( .in(\mat_add/r102/B_AS [4]), .out(
        \mat_mul/mult_37_G2_G1_G1/B_not [4]) );
  inv \mat_mul/mult_37_G2_G1_G1/AN1_3_0  ( .in(\mat_add/r102/B_AS [3]), .out(
        \mat_mul/mult_37_G2_G1_G1/B_not [3]) );
  inv \mat_mul/mult_37_G2_G1_G1/AN1_2_0  ( .in(\mat_add/r102/B_AS [2]), .out(
        \mat_mul/mult_37_G2_G1_G1/B_not [2]) );
  inv \mat_mul/mult_37_G2_G1_G1/AN1_1_0  ( .in(\mat_add/r102/B_AS [1]), .out(
        \mat_mul/mult_37_G2_G1_G1/B_not [1]) );
  inv \mat_mul/mult_37_G2_G1_G1/AN1_0_0  ( .in(\mat_add/r102/B_AS [0]), .out(
        \mat_mul/mult_37_G2_G1_G1/B_notx[0] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN3_7_0  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [7]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[7][0] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_6_1  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [6]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[6][1] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_6_0_0  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [6]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[6][0] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_5_2  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [5]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[5][2] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_5_1  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [5]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[5][1] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_5_0_0  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [5]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[5][0] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_4_3  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [4]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [3]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[4][3] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_4_2  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [4]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[4][2] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_4_1  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [4]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[4][1] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_4_0_0  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [4]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[4][0] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_3_4  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [3]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [4]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[3][4] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_3_3  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [3]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [3]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[3][3] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_3_2  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [3]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[3][2] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_3_1  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [3]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[3][1] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_3_0_0  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [3]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[3][0] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_2_5  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [2]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [5]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[2][5] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_2_4  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [2]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [4]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[2][4] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_2_3  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [2]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [3]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[2][3] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_2_2  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [2]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[2][2] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_2_1  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [2]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[2][1] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_2_0_0  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [2]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[2][0] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_1_6  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [1]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [6]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[1][6] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_1_5  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [1]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [5]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[1][5] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_1_4  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [1]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [4]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[1][4] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_1_3  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [1]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [3]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[1][3] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_1_2  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [1]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[1][2] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_1_1  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [1]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[1][1] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_1_0_0  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_not [1]), .b(
        \mat_mul/mult_37_G2_G1_G1/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[1][0] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN2_0_7  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [7]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[0][7] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_0_6  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [6]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[0][6] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_0_5  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [5]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[0][5] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_0_4  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [4]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[0][4] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_0_3  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [3]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[0][3] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_0_2  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[0][2] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_0_1  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G1_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1_G1/ab[0][1] ) );
  nor2 \mat_mul/mult_37_G2_G1_G1/AN1_0_0_0  ( .a(
        \mat_mul/mult_37_G2_G1_G1/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G1_G1/B_notx[0] ), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[0] ) );
  inv \mat_mul/mult_37_G2_G1/AN1_7  ( .in(A[31]), .out(
        \mat_mul/mult_37_G2_G1/A_not [7]) );
  inv \mat_mul/mult_37_G2_G1/AN1_6  ( .in(A[30]), .out(
        \mat_mul/mult_37_G2_G1/A_not [6]) );
  inv \mat_mul/mult_37_G2_G1/AN1_5  ( .in(A[29]), .out(
        \mat_mul/mult_37_G2_G1/A_not [5]) );
  inv \mat_mul/mult_37_G2_G1/AN1_4  ( .in(A[28]), .out(
        \mat_mul/mult_37_G2_G1/A_not [4]) );
  inv \mat_mul/mult_37_G2_G1/AN1_3  ( .in(A[27]), .out(
        \mat_mul/mult_37_G2_G1/A_not [3]) );
  inv \mat_mul/mult_37_G2_G1/AN1_2  ( .in(A[26]), .out(
        \mat_mul/mult_37_G2_G1/A_not [2]) );
  inv \mat_mul/mult_37_G2_G1/AN1_1  ( .in(A[25]), .out(
        \mat_mul/mult_37_G2_G1/A_not [1]) );
  inv \mat_mul/mult_37_G2_G1/AN1_0  ( .in(A[24]), .out(
        \mat_mul/mult_37_G2_G1/A_notx[0] ) );
  inv \mat_mul/mult_37_G2_G1/AN1_7_0  ( .in(\mat_add/r98/B_AS [7]), .out(
        \mat_mul/mult_37_G2_G1/B_not [7]) );
  inv \mat_mul/mult_37_G2_G1/AN1_6_0  ( .in(\mat_add/r98/B_AS [6]), .out(
        \mat_mul/mult_37_G2_G1/B_not [6]) );
  inv \mat_mul/mult_37_G2_G1/AN1_5_0  ( .in(\mat_add/r98/B_AS [5]), .out(
        \mat_mul/mult_37_G2_G1/B_not [5]) );
  inv \mat_mul/mult_37_G2_G1/AN1_4_0  ( .in(\mat_add/r98/B_AS [4]), .out(
        \mat_mul/mult_37_G2_G1/B_not [4]) );
  inv \mat_mul/mult_37_G2_G1/AN1_3_0  ( .in(\mat_add/r98/B_AS [3]), .out(
        \mat_mul/mult_37_G2_G1/B_not [3]) );
  inv \mat_mul/mult_37_G2_G1/AN1_2_0  ( .in(\mat_add/r98/B_AS [2]), .out(
        \mat_mul/mult_37_G2_G1/B_not [2]) );
  inv \mat_mul/mult_37_G2_G1/AN1_1_0  ( .in(\mat_add/r98/B_AS [1]), .out(
        \mat_mul/mult_37_G2_G1/B_not [1]) );
  inv \mat_mul/mult_37_G2_G1/AN1_0_0  ( .in(\mat_add/r98/B_AS [0]), .out(
        \mat_mul/mult_37_G2_G1/B_notx[0] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN3_7_0  ( .a(\mat_mul/mult_37_G2_G1/A_not [7]), 
        .b(\mat_mul/mult_37_G2_G1/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G1/ab[7][0] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_6_1  ( .a(\mat_mul/mult_37_G2_G1/A_not [6]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1/ab[6][1] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_6_0_0  ( .a(\mat_mul/mult_37_G2_G1/A_not [6]), .b(\mat_mul/mult_37_G2_G1/B_notx[0] ), .out(\mat_mul/mult_37_G2_G1/ab[6][0] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_5_2  ( .a(\mat_mul/mult_37_G2_G1/A_not [5]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1/ab[5][2] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_5_1  ( .a(\mat_mul/mult_37_G2_G1/A_not [5]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1/ab[5][1] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_5_0_0  ( .a(\mat_mul/mult_37_G2_G1/A_not [5]), .b(\mat_mul/mult_37_G2_G1/B_notx[0] ), .out(\mat_mul/mult_37_G2_G1/ab[5][0] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_4_3  ( .a(\mat_mul/mult_37_G2_G1/A_not [4]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [3]), .out(
        \mat_mul/mult_37_G2_G1/ab[4][3] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_4_2  ( .a(\mat_mul/mult_37_G2_G1/A_not [4]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1/ab[4][2] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_4_1  ( .a(\mat_mul/mult_37_G2_G1/A_not [4]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1/ab[4][1] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_4_0_0  ( .a(\mat_mul/mult_37_G2_G1/A_not [4]), .b(\mat_mul/mult_37_G2_G1/B_notx[0] ), .out(\mat_mul/mult_37_G2_G1/ab[4][0] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_3_4  ( .a(\mat_mul/mult_37_G2_G1/A_not [3]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [4]), .out(
        \mat_mul/mult_37_G2_G1/ab[3][4] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_3_3  ( .a(\mat_mul/mult_37_G2_G1/A_not [3]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [3]), .out(
        \mat_mul/mult_37_G2_G1/ab[3][3] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_3_2  ( .a(\mat_mul/mult_37_G2_G1/A_not [3]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1/ab[3][2] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_3_1  ( .a(\mat_mul/mult_37_G2_G1/A_not [3]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1/ab[3][1] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_3_0_0  ( .a(\mat_mul/mult_37_G2_G1/A_not [3]), .b(\mat_mul/mult_37_G2_G1/B_notx[0] ), .out(\mat_mul/mult_37_G2_G1/ab[3][0] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_2_5  ( .a(\mat_mul/mult_37_G2_G1/A_not [2]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [5]), .out(
        \mat_mul/mult_37_G2_G1/ab[2][5] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_2_4  ( .a(\mat_mul/mult_37_G2_G1/A_not [2]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [4]), .out(
        \mat_mul/mult_37_G2_G1/ab[2][4] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_2_3  ( .a(\mat_mul/mult_37_G2_G1/A_not [2]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [3]), .out(
        \mat_mul/mult_37_G2_G1/ab[2][3] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_2_2  ( .a(\mat_mul/mult_37_G2_G1/A_not [2]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1/ab[2][2] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_2_1  ( .a(\mat_mul/mult_37_G2_G1/A_not [2]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1/ab[2][1] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_2_0_0  ( .a(\mat_mul/mult_37_G2_G1/A_not [2]), .b(\mat_mul/mult_37_G2_G1/B_notx[0] ), .out(\mat_mul/mult_37_G2_G1/ab[2][0] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_1_6  ( .a(\mat_mul/mult_37_G2_G1/A_not [1]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [6]), .out(
        \mat_mul/mult_37_G2_G1/ab[1][6] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_1_5  ( .a(\mat_mul/mult_37_G2_G1/A_not [1]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [5]), .out(
        \mat_mul/mult_37_G2_G1/ab[1][5] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_1_4  ( .a(\mat_mul/mult_37_G2_G1/A_not [1]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [4]), .out(
        \mat_mul/mult_37_G2_G1/ab[1][4] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_1_3  ( .a(\mat_mul/mult_37_G2_G1/A_not [1]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [3]), .out(
        \mat_mul/mult_37_G2_G1/ab[1][3] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_1_2  ( .a(\mat_mul/mult_37_G2_G1/A_not [1]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1/ab[1][2] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_1_1  ( .a(\mat_mul/mult_37_G2_G1/A_not [1]), 
        .b(\mat_mul/mult_37_G2_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1/ab[1][1] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_1_0_0  ( .a(\mat_mul/mult_37_G2_G1/A_not [1]), .b(\mat_mul/mult_37_G2_G1/B_notx[0] ), .out(\mat_mul/mult_37_G2_G1/ab[1][0] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN2_0_7  ( .a(\mat_mul/mult_37_G2_G1/A_notx[0] ), 
        .b(\mat_mul/mult_37_G2_G1/B_not [7]), .out(
        \mat_mul/mult_37_G2_G1/ab[0][7] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_0_6  ( .a(\mat_mul/mult_37_G2_G1/A_notx[0] ), 
        .b(\mat_mul/mult_37_G2_G1/B_not [6]), .out(
        \mat_mul/mult_37_G2_G1/ab[0][6] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_0_5  ( .a(\mat_mul/mult_37_G2_G1/A_notx[0] ), 
        .b(\mat_mul/mult_37_G2_G1/B_not [5]), .out(
        \mat_mul/mult_37_G2_G1/ab[0][5] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_0_4  ( .a(\mat_mul/mult_37_G2_G1/A_notx[0] ), 
        .b(\mat_mul/mult_37_G2_G1/B_not [4]), .out(
        \mat_mul/mult_37_G2_G1/ab[0][4] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_0_3  ( .a(\mat_mul/mult_37_G2_G1/A_notx[0] ), 
        .b(\mat_mul/mult_37_G2_G1/B_not [3]), .out(
        \mat_mul/mult_37_G2_G1/ab[0][3] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_0_2  ( .a(\mat_mul/mult_37_G2_G1/A_notx[0] ), 
        .b(\mat_mul/mult_37_G2_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1/ab[0][2] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_0_1  ( .a(\mat_mul/mult_37_G2_G1/A_notx[0] ), 
        .b(\mat_mul/mult_37_G2_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1/ab[0][1] ) );
  nor2 \mat_mul/mult_37_G2_G1/AN1_0_0_0  ( .a(
        \mat_mul/mult_37_G2_G1/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G1/B_notx[0] ), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[0] ) );
  inv \mat_mul/mult_37_G2_G2_G1/AN1_7  ( .in(A[23]), .out(
        \mat_mul/mult_37_G2_G2_G1/A_not [7]) );
  inv \mat_mul/mult_37_G2_G2_G1/AN1_6  ( .in(A[22]), .out(
        \mat_mul/mult_37_G2_G2_G1/A_not [6]) );
  inv \mat_mul/mult_37_G2_G2_G1/AN1_5  ( .in(A[21]), .out(
        \mat_mul/mult_37_G2_G2_G1/A_not [5]) );
  inv \mat_mul/mult_37_G2_G2_G1/AN1_4  ( .in(A[20]), .out(
        \mat_mul/mult_37_G2_G2_G1/A_not [4]) );
  inv \mat_mul/mult_37_G2_G2_G1/AN1_3  ( .in(A[19]), .out(
        \mat_mul/mult_37_G2_G2_G1/A_not [3]) );
  inv \mat_mul/mult_37_G2_G2_G1/AN1_2  ( .in(A[18]), .out(
        \mat_mul/mult_37_G2_G2_G1/A_not [2]) );
  inv \mat_mul/mult_37_G2_G2_G1/AN1_1  ( .in(A[17]), .out(
        \mat_mul/mult_37_G2_G2_G1/A_not [1]) );
  inv \mat_mul/mult_37_G2_G2_G1/AN1_0  ( .in(A[16]), .out(
        \mat_mul/mult_37_G2_G2_G1/A_notx[0] ) );
  inv \mat_mul/mult_37_G2_G2_G1/AN1_7_0  ( .in(\mat_add/r106/B_AS [7]), .out(
        \mat_mul/mult_37_G2_G2_G1/B_not [7]) );
  inv \mat_mul/mult_37_G2_G2_G1/AN1_6_0  ( .in(\mat_add/r106/B_AS [6]), .out(
        \mat_mul/mult_37_G2_G2_G1/B_not [6]) );
  inv \mat_mul/mult_37_G2_G2_G1/AN1_5_0  ( .in(\mat_add/r106/B_AS [5]), .out(
        \mat_mul/mult_37_G2_G2_G1/B_not [5]) );
  inv \mat_mul/mult_37_G2_G2_G1/AN1_4_0  ( .in(\mat_add/r106/B_AS [4]), .out(
        \mat_mul/mult_37_G2_G2_G1/B_not [4]) );
  inv \mat_mul/mult_37_G2_G2_G1/AN1_3_0  ( .in(\mat_add/r106/B_AS [3]), .out(
        \mat_mul/mult_37_G2_G2_G1/B_not [3]) );
  inv \mat_mul/mult_37_G2_G2_G1/AN1_2_0  ( .in(\mat_add/r106/B_AS [2]), .out(
        \mat_mul/mult_37_G2_G2_G1/B_not [2]) );
  inv \mat_mul/mult_37_G2_G2_G1/AN1_1_0  ( .in(\mat_add/r106/B_AS [1]), .out(
        \mat_mul/mult_37_G2_G2_G1/B_not [1]) );
  inv \mat_mul/mult_37_G2_G2_G1/AN1_0_0  ( .in(\mat_add/r106/B_AS [0]), .out(
        \mat_mul/mult_37_G2_G2_G1/B_notx[0] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN3_7_0  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [7]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[7][0] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_6_1  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [6]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[6][1] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_6_0_0  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [6]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[6][0] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_5_2  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [5]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[5][2] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_5_1  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [5]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[5][1] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_5_0_0  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [5]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[5][0] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_4_3  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [4]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [3]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[4][3] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_4_2  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [4]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[4][2] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_4_1  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [4]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[4][1] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_4_0_0  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [4]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[4][0] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_3_4  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [3]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [4]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[3][4] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_3_3  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [3]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [3]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[3][3] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_3_2  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [3]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[3][2] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_3_1  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [3]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[3][1] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_3_0_0  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [3]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[3][0] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_2_5  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [2]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [5]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[2][5] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_2_4  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [2]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [4]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[2][4] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_2_3  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [2]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [3]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[2][3] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_2_2  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [2]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[2][2] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_2_1  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [2]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[2][1] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_2_0_0  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [2]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[2][0] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_1_6  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [1]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [6]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[1][6] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_1_5  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [1]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [5]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[1][5] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_1_4  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [1]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [4]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[1][4] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_1_3  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [1]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [3]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[1][3] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_1_2  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [1]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[1][2] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_1_1  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [1]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[1][1] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_1_0_0  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_not [1]), .b(
        \mat_mul/mult_37_G2_G2_G1/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[1][0] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN2_0_7  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [7]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[0][7] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_0_6  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [6]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[0][6] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_0_5  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [5]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[0][5] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_0_4  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [4]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[0][4] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_0_3  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [3]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[0][3] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_0_2  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[0][2] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_0_1  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G2_G1/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2_G1/ab[0][1] ) );
  nor2 \mat_mul/mult_37_G2_G2_G1/AN1_0_0_0  ( .a(
        \mat_mul/mult_37_G2_G2_G1/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G2_G1/B_notx[0] ), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[0] ) );
  inv \mat_mul/mult_37_G2/AN1_7  ( .in(A[15]), .out(
        \mat_mul/mult_37_G2/A_not [7]) );
  inv \mat_mul/mult_37_G2/AN1_6  ( .in(A[14]), .out(
        \mat_mul/mult_37_G2/A_not [6]) );
  inv \mat_mul/mult_37_G2/AN1_5  ( .in(A[13]), .out(
        \mat_mul/mult_37_G2/A_not [5]) );
  inv \mat_mul/mult_37_G2/AN1_4  ( .in(A[12]), .out(
        \mat_mul/mult_37_G2/A_not [4]) );
  inv \mat_mul/mult_37_G2/AN1_3  ( .in(A[11]), .out(
        \mat_mul/mult_37_G2/A_not [3]) );
  inv \mat_mul/mult_37_G2/AN1_2  ( .in(A[10]), .out(
        \mat_mul/mult_37_G2/A_not [2]) );
  inv \mat_mul/mult_37_G2/AN1_1  ( .in(A[9]), .out(
        \mat_mul/mult_37_G2/A_not [1]) );
  inv \mat_mul/mult_37_G2/AN1_0  ( .in(A[8]), .out(
        \mat_mul/mult_37_G2/A_notx[0] ) );
  inv \mat_mul/mult_37_G2/AN1_7_0  ( .in(\mat_add/r94/B_AS [7]), .out(
        \mat_mul/mult_37_G2/B_not [7]) );
  inv \mat_mul/mult_37_G2/AN1_6_0  ( .in(\mat_add/r94/B_AS [6]), .out(
        \mat_mul/mult_37_G2/B_not [6]) );
  inv \mat_mul/mult_37_G2/AN1_5_0  ( .in(\mat_add/r94/B_AS [5]), .out(
        \mat_mul/mult_37_G2/B_not [5]) );
  inv \mat_mul/mult_37_G2/AN1_4_0  ( .in(\mat_add/r94/B_AS [4]), .out(
        \mat_mul/mult_37_G2/B_not [4]) );
  inv \mat_mul/mult_37_G2/AN1_3_0  ( .in(\mat_add/r94/B_AS [3]), .out(
        \mat_mul/mult_37_G2/B_not [3]) );
  inv \mat_mul/mult_37_G2/AN1_2_0  ( .in(\mat_add/r94/B_AS [2]), .out(
        \mat_mul/mult_37_G2/B_not [2]) );
  inv \mat_mul/mult_37_G2/AN1_1_0  ( .in(\mat_add/r94/B_AS [1]), .out(
        \mat_mul/mult_37_G2/B_not [1]) );
  inv \mat_mul/mult_37_G2/AN1_0_0  ( .in(\mat_add/r94/B_AS [0]), .out(
        \mat_mul/mult_37_G2/B_notx[0] ) );
  nor2 \mat_mul/mult_37_G2/AN3_7_0  ( .a(\mat_mul/mult_37_G2/A_not [7]), .b(
        \mat_mul/mult_37_G2/B_notx[0] ), .out(\mat_mul/mult_37_G2/ab[7][0] )
         );
  nor2 \mat_mul/mult_37_G2/AN1_6_1  ( .a(\mat_mul/mult_37_G2/A_not [6]), .b(
        \mat_mul/mult_37_G2/B_not [1]), .out(\mat_mul/mult_37_G2/ab[6][1] ) );
  nor2 \mat_mul/mult_37_G2/AN1_6_0_0  ( .a(\mat_mul/mult_37_G2/A_not [6]), .b(
        \mat_mul/mult_37_G2/B_notx[0] ), .out(\mat_mul/mult_37_G2/ab[6][0] )
         );
  nor2 \mat_mul/mult_37_G2/AN1_5_2  ( .a(\mat_mul/mult_37_G2/A_not [5]), .b(
        \mat_mul/mult_37_G2/B_not [2]), .out(\mat_mul/mult_37_G2/ab[5][2] ) );
  nor2 \mat_mul/mult_37_G2/AN1_5_1  ( .a(\mat_mul/mult_37_G2/A_not [5]), .b(
        \mat_mul/mult_37_G2/B_not [1]), .out(\mat_mul/mult_37_G2/ab[5][1] ) );
  nor2 \mat_mul/mult_37_G2/AN1_5_0_0  ( .a(\mat_mul/mult_37_G2/A_not [5]), .b(
        \mat_mul/mult_37_G2/B_notx[0] ), .out(\mat_mul/mult_37_G2/ab[5][0] )
         );
  nor2 \mat_mul/mult_37_G2/AN1_4_3  ( .a(\mat_mul/mult_37_G2/A_not [4]), .b(
        \mat_mul/mult_37_G2/B_not [3]), .out(\mat_mul/mult_37_G2/ab[4][3] ) );
  nor2 \mat_mul/mult_37_G2/AN1_4_2  ( .a(\mat_mul/mult_37_G2/A_not [4]), .b(
        \mat_mul/mult_37_G2/B_not [2]), .out(\mat_mul/mult_37_G2/ab[4][2] ) );
  nor2 \mat_mul/mult_37_G2/AN1_4_1  ( .a(\mat_mul/mult_37_G2/A_not [4]), .b(
        \mat_mul/mult_37_G2/B_not [1]), .out(\mat_mul/mult_37_G2/ab[4][1] ) );
  nor2 \mat_mul/mult_37_G2/AN1_4_0_0  ( .a(\mat_mul/mult_37_G2/A_not [4]), .b(
        \mat_mul/mult_37_G2/B_notx[0] ), .out(\mat_mul/mult_37_G2/ab[4][0] )
         );
  nor2 \mat_mul/mult_37_G2/AN1_3_4  ( .a(\mat_mul/mult_37_G2/A_not [3]), .b(
        \mat_mul/mult_37_G2/B_not [4]), .out(\mat_mul/mult_37_G2/ab[3][4] ) );
  nor2 \mat_mul/mult_37_G2/AN1_3_3  ( .a(\mat_mul/mult_37_G2/A_not [3]), .b(
        \mat_mul/mult_37_G2/B_not [3]), .out(\mat_mul/mult_37_G2/ab[3][3] ) );
  nor2 \mat_mul/mult_37_G2/AN1_3_2  ( .a(\mat_mul/mult_37_G2/A_not [3]), .b(
        \mat_mul/mult_37_G2/B_not [2]), .out(\mat_mul/mult_37_G2/ab[3][2] ) );
  nor2 \mat_mul/mult_37_G2/AN1_3_1  ( .a(\mat_mul/mult_37_G2/A_not [3]), .b(
        \mat_mul/mult_37_G2/B_not [1]), .out(\mat_mul/mult_37_G2/ab[3][1] ) );
  nor2 \mat_mul/mult_37_G2/AN1_3_0_0  ( .a(\mat_mul/mult_37_G2/A_not [3]), .b(
        \mat_mul/mult_37_G2/B_notx[0] ), .out(\mat_mul/mult_37_G2/ab[3][0] )
         );
  nor2 \mat_mul/mult_37_G2/AN1_2_5  ( .a(\mat_mul/mult_37_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2/B_not [5]), .out(\mat_mul/mult_37_G2/ab[2][5] ) );
  nor2 \mat_mul/mult_37_G2/AN1_2_4  ( .a(\mat_mul/mult_37_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2/B_not [4]), .out(\mat_mul/mult_37_G2/ab[2][4] ) );
  nor2 \mat_mul/mult_37_G2/AN1_2_3  ( .a(\mat_mul/mult_37_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2/B_not [3]), .out(\mat_mul/mult_37_G2/ab[2][3] ) );
  nor2 \mat_mul/mult_37_G2/AN1_2_2  ( .a(\mat_mul/mult_37_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2/B_not [2]), .out(\mat_mul/mult_37_G2/ab[2][2] ) );
  nor2 \mat_mul/mult_37_G2/AN1_2_1  ( .a(\mat_mul/mult_37_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2/B_not [1]), .out(\mat_mul/mult_37_G2/ab[2][1] ) );
  nor2 \mat_mul/mult_37_G2/AN1_2_0_0  ( .a(\mat_mul/mult_37_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2/B_notx[0] ), .out(\mat_mul/mult_37_G2/ab[2][0] )
         );
  nor2 \mat_mul/mult_37_G2/AN1_1_6  ( .a(\mat_mul/mult_37_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2/B_not [6]), .out(\mat_mul/mult_37_G2/ab[1][6] ) );
  nor2 \mat_mul/mult_37_G2/AN1_1_5  ( .a(\mat_mul/mult_37_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2/B_not [5]), .out(\mat_mul/mult_37_G2/ab[1][5] ) );
  nor2 \mat_mul/mult_37_G2/AN1_1_4  ( .a(\mat_mul/mult_37_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2/B_not [4]), .out(\mat_mul/mult_37_G2/ab[1][4] ) );
  nor2 \mat_mul/mult_37_G2/AN1_1_3  ( .a(\mat_mul/mult_37_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2/B_not [3]), .out(\mat_mul/mult_37_G2/ab[1][3] ) );
  nor2 \mat_mul/mult_37_G2/AN1_1_2  ( .a(\mat_mul/mult_37_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2/B_not [2]), .out(\mat_mul/mult_37_G2/ab[1][2] ) );
  nor2 \mat_mul/mult_37_G2/AN1_1_1  ( .a(\mat_mul/mult_37_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2/B_not [1]), .out(\mat_mul/mult_37_G2/ab[1][1] ) );
  nor2 \mat_mul/mult_37_G2/AN1_1_0_0  ( .a(\mat_mul/mult_37_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2/B_notx[0] ), .out(\mat_mul/mult_37_G2/ab[1][0] )
         );
  nor2 \mat_mul/mult_37_G2/AN2_0_7  ( .a(\mat_mul/mult_37_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2/B_not [7]), .out(\mat_mul/mult_37_G2/ab[0][7] ) );
  nor2 \mat_mul/mult_37_G2/AN1_0_6  ( .a(\mat_mul/mult_37_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2/B_not [6]), .out(\mat_mul/mult_37_G2/ab[0][6] ) );
  nor2 \mat_mul/mult_37_G2/AN1_0_5  ( .a(\mat_mul/mult_37_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2/B_not [5]), .out(\mat_mul/mult_37_G2/ab[0][5] ) );
  nor2 \mat_mul/mult_37_G2/AN1_0_4  ( .a(\mat_mul/mult_37_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2/B_not [4]), .out(\mat_mul/mult_37_G2/ab[0][4] ) );
  nor2 \mat_mul/mult_37_G2/AN1_0_3  ( .a(\mat_mul/mult_37_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2/B_not [3]), .out(\mat_mul/mult_37_G2/ab[0][3] ) );
  nor2 \mat_mul/mult_37_G2/AN1_0_2  ( .a(\mat_mul/mult_37_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2/B_not [2]), .out(\mat_mul/mult_37_G2/ab[0][2] ) );
  nor2 \mat_mul/mult_37_G2/AN1_0_1  ( .a(\mat_mul/mult_37_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2/B_not [1]), .out(\mat_mul/mult_37_G2/ab[0][1] ) );
  nor2 \mat_mul/mult_37_G2/AN1_0_0_0  ( .a(\mat_mul/mult_37_G2/A_notx[0] ), 
        .b(\mat_mul/mult_37_G2/B_notx[0] ), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[0] ) );
  inv \mat_mul/mult_37_G2_G1_G2/AN1_7  ( .in(A[7]), .out(
        \mat_mul/mult_37_G2_G1_G2/A_not [7]) );
  inv \mat_mul/mult_37_G2_G1_G2/AN1_6  ( .in(A[6]), .out(
        \mat_mul/mult_37_G2_G1_G2/A_not [6]) );
  inv \mat_mul/mult_37_G2_G1_G2/AN1_5  ( .in(A[5]), .out(
        \mat_mul/mult_37_G2_G1_G2/A_not [5]) );
  inv \mat_mul/mult_37_G2_G1_G2/AN1_4  ( .in(A[4]), .out(
        \mat_mul/mult_37_G2_G1_G2/A_not [4]) );
  inv \mat_mul/mult_37_G2_G1_G2/AN1_3  ( .in(A[3]), .out(
        \mat_mul/mult_37_G2_G1_G2/A_not [3]) );
  inv \mat_mul/mult_37_G2_G1_G2/AN1_2  ( .in(A[2]), .out(
        \mat_mul/mult_37_G2_G1_G2/A_not [2]) );
  inv \mat_mul/mult_37_G2_G1_G2/AN1_1  ( .in(A[1]), .out(
        \mat_mul/mult_37_G2_G1_G2/A_not [1]) );
  inv \mat_mul/mult_37_G2_G1_G2/AN1_0  ( .in(A[0]), .out(
        \mat_mul/mult_37_G2_G1_G2/A_notx[0] ) );
  inv \mat_mul/mult_37_G2_G1_G2/AN1_7_0  ( .in(\mat_add/r102/B_AS [7]), .out(
        \mat_mul/mult_37_G2_G1_G2/B_not [7]) );
  inv \mat_mul/mult_37_G2_G1_G2/AN1_6_0  ( .in(\mat_add/r102/B_AS [6]), .out(
        \mat_mul/mult_37_G2_G1_G2/B_not [6]) );
  inv \mat_mul/mult_37_G2_G1_G2/AN1_5_0  ( .in(\mat_add/r102/B_AS [5]), .out(
        \mat_mul/mult_37_G2_G1_G2/B_not [5]) );
  inv \mat_mul/mult_37_G2_G1_G2/AN1_4_0  ( .in(\mat_add/r102/B_AS [4]), .out(
        \mat_mul/mult_37_G2_G1_G2/B_not [4]) );
  inv \mat_mul/mult_37_G2_G1_G2/AN1_3_0  ( .in(\mat_add/r102/B_AS [3]), .out(
        \mat_mul/mult_37_G2_G1_G2/B_not [3]) );
  inv \mat_mul/mult_37_G2_G1_G2/AN1_2_0  ( .in(\mat_add/r102/B_AS [2]), .out(
        \mat_mul/mult_37_G2_G1_G2/B_not [2]) );
  inv \mat_mul/mult_37_G2_G1_G2/AN1_1_0  ( .in(\mat_add/r102/B_AS [1]), .out(
        \mat_mul/mult_37_G2_G1_G2/B_not [1]) );
  inv \mat_mul/mult_37_G2_G1_G2/AN1_0_0  ( .in(\mat_add/r102/B_AS [0]), .out(
        \mat_mul/mult_37_G2_G1_G2/B_notx[0] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN3_7_0  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [7]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[7][0] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_6_1  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [6]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[6][1] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_6_0_0  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [6]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[6][0] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_5_2  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [5]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[5][2] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_5_1  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [5]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[5][1] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_5_0_0  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [5]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[5][0] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_4_3  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [4]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [3]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[4][3] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_4_2  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [4]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[4][2] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_4_1  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [4]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[4][1] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_4_0_0  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [4]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[4][0] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_3_4  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [3]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [4]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[3][4] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_3_3  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [3]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [3]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[3][3] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_3_2  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [3]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[3][2] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_3_1  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [3]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[3][1] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_3_0_0  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [3]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[3][0] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_2_5  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [5]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[2][5] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_2_4  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [4]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[2][4] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_2_3  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [3]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[2][3] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_2_2  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[2][2] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_2_1  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[2][1] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_2_0_0  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[2][0] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_1_6  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [6]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[1][6] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_1_5  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [5]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[1][5] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_1_4  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [4]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[1][4] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_1_3  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [3]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[1][3] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_1_2  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[1][2] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_1_1  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[1][1] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_1_0_0  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2_G1_G2/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[1][0] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN2_0_7  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [7]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[0][7] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_0_6  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [6]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[0][6] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_0_5  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [5]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[0][5] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_0_4  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [4]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[0][4] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_0_3  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [3]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[0][3] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_0_2  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[0][2] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_0_1  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G1_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G1_G2/ab[0][1] ) );
  nor2 \mat_mul/mult_37_G2_G1_G2/AN1_0_0_0  ( .a(
        \mat_mul/mult_37_G2_G1_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G1_G2/B_notx[0] ), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[0] ) );
  inv \mat_mul/mult_37_G2_G2/AN1_7  ( .in(A[15]), .out(
        \mat_mul/mult_37_G2_G2/A_not [7]) );
  inv \mat_mul/mult_37_G2_G2/AN1_6  ( .in(A[14]), .out(
        \mat_mul/mult_37_G2_G2/A_not [6]) );
  inv \mat_mul/mult_37_G2_G2/AN1_5  ( .in(A[13]), .out(
        \mat_mul/mult_37_G2_G2/A_not [5]) );
  inv \mat_mul/mult_37_G2_G2/AN1_4  ( .in(A[12]), .out(
        \mat_mul/mult_37_G2_G2/A_not [4]) );
  inv \mat_mul/mult_37_G2_G2/AN1_3  ( .in(A[11]), .out(
        \mat_mul/mult_37_G2_G2/A_not [3]) );
  inv \mat_mul/mult_37_G2_G2/AN1_2  ( .in(A[10]), .out(
        \mat_mul/mult_37_G2_G2/A_not [2]) );
  inv \mat_mul/mult_37_G2_G2/AN1_1  ( .in(A[9]), .out(
        \mat_mul/mult_37_G2_G2/A_not [1]) );
  inv \mat_mul/mult_37_G2_G2/AN1_0  ( .in(A[8]), .out(
        \mat_mul/mult_37_G2_G2/A_notx[0] ) );
  inv \mat_mul/mult_37_G2_G2/AN1_7_0  ( .in(\mat_add/r98/B_AS [7]), .out(
        \mat_mul/mult_37_G2_G2/B_not [7]) );
  inv \mat_mul/mult_37_G2_G2/AN1_6_0  ( .in(\mat_add/r98/B_AS [6]), .out(
        \mat_mul/mult_37_G2_G2/B_not [6]) );
  inv \mat_mul/mult_37_G2_G2/AN1_5_0  ( .in(\mat_add/r98/B_AS [5]), .out(
        \mat_mul/mult_37_G2_G2/B_not [5]) );
  inv \mat_mul/mult_37_G2_G2/AN1_4_0  ( .in(\mat_add/r98/B_AS [4]), .out(
        \mat_mul/mult_37_G2_G2/B_not [4]) );
  inv \mat_mul/mult_37_G2_G2/AN1_3_0  ( .in(\mat_add/r98/B_AS [3]), .out(
        \mat_mul/mult_37_G2_G2/B_not [3]) );
  inv \mat_mul/mult_37_G2_G2/AN1_2_0  ( .in(\mat_add/r98/B_AS [2]), .out(
        \mat_mul/mult_37_G2_G2/B_not [2]) );
  inv \mat_mul/mult_37_G2_G2/AN1_1_0  ( .in(\mat_add/r98/B_AS [1]), .out(
        \mat_mul/mult_37_G2_G2/B_not [1]) );
  inv \mat_mul/mult_37_G2_G2/AN1_0_0  ( .in(\mat_add/r98/B_AS [0]), .out(
        \mat_mul/mult_37_G2_G2/B_notx[0] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN3_7_0  ( .a(\mat_mul/mult_37_G2_G2/A_not [7]), 
        .b(\mat_mul/mult_37_G2_G2/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G2/ab[7][0] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_6_1  ( .a(\mat_mul/mult_37_G2_G2/A_not [6]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2/ab[6][1] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_6_0_0  ( .a(\mat_mul/mult_37_G2_G2/A_not [6]), .b(\mat_mul/mult_37_G2_G2/B_notx[0] ), .out(\mat_mul/mult_37_G2_G2/ab[6][0] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_5_2  ( .a(\mat_mul/mult_37_G2_G2/A_not [5]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2/ab[5][2] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_5_1  ( .a(\mat_mul/mult_37_G2_G2/A_not [5]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2/ab[5][1] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_5_0_0  ( .a(\mat_mul/mult_37_G2_G2/A_not [5]), .b(\mat_mul/mult_37_G2_G2/B_notx[0] ), .out(\mat_mul/mult_37_G2_G2/ab[5][0] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_4_3  ( .a(\mat_mul/mult_37_G2_G2/A_not [4]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [3]), .out(
        \mat_mul/mult_37_G2_G2/ab[4][3] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_4_2  ( .a(\mat_mul/mult_37_G2_G2/A_not [4]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2/ab[4][2] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_4_1  ( .a(\mat_mul/mult_37_G2_G2/A_not [4]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2/ab[4][1] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_4_0_0  ( .a(\mat_mul/mult_37_G2_G2/A_not [4]), .b(\mat_mul/mult_37_G2_G2/B_notx[0] ), .out(\mat_mul/mult_37_G2_G2/ab[4][0] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_3_4  ( .a(\mat_mul/mult_37_G2_G2/A_not [3]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [4]), .out(
        \mat_mul/mult_37_G2_G2/ab[3][4] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_3_3  ( .a(\mat_mul/mult_37_G2_G2/A_not [3]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [3]), .out(
        \mat_mul/mult_37_G2_G2/ab[3][3] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_3_2  ( .a(\mat_mul/mult_37_G2_G2/A_not [3]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2/ab[3][2] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_3_1  ( .a(\mat_mul/mult_37_G2_G2/A_not [3]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2/ab[3][1] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_3_0_0  ( .a(\mat_mul/mult_37_G2_G2/A_not [3]), .b(\mat_mul/mult_37_G2_G2/B_notx[0] ), .out(\mat_mul/mult_37_G2_G2/ab[3][0] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_2_5  ( .a(\mat_mul/mult_37_G2_G2/A_not [2]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [5]), .out(
        \mat_mul/mult_37_G2_G2/ab[2][5] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_2_4  ( .a(\mat_mul/mult_37_G2_G2/A_not [2]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [4]), .out(
        \mat_mul/mult_37_G2_G2/ab[2][4] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_2_3  ( .a(\mat_mul/mult_37_G2_G2/A_not [2]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [3]), .out(
        \mat_mul/mult_37_G2_G2/ab[2][3] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_2_2  ( .a(\mat_mul/mult_37_G2_G2/A_not [2]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2/ab[2][2] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_2_1  ( .a(\mat_mul/mult_37_G2_G2/A_not [2]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2/ab[2][1] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_2_0_0  ( .a(\mat_mul/mult_37_G2_G2/A_not [2]), .b(\mat_mul/mult_37_G2_G2/B_notx[0] ), .out(\mat_mul/mult_37_G2_G2/ab[2][0] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_1_6  ( .a(\mat_mul/mult_37_G2_G2/A_not [1]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [6]), .out(
        \mat_mul/mult_37_G2_G2/ab[1][6] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_1_5  ( .a(\mat_mul/mult_37_G2_G2/A_not [1]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [5]), .out(
        \mat_mul/mult_37_G2_G2/ab[1][5] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_1_4  ( .a(\mat_mul/mult_37_G2_G2/A_not [1]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [4]), .out(
        \mat_mul/mult_37_G2_G2/ab[1][4] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_1_3  ( .a(\mat_mul/mult_37_G2_G2/A_not [1]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [3]), .out(
        \mat_mul/mult_37_G2_G2/ab[1][3] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_1_2  ( .a(\mat_mul/mult_37_G2_G2/A_not [1]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2/ab[1][2] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_1_1  ( .a(\mat_mul/mult_37_G2_G2/A_not [1]), 
        .b(\mat_mul/mult_37_G2_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2/ab[1][1] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_1_0_0  ( .a(\mat_mul/mult_37_G2_G2/A_not [1]), .b(\mat_mul/mult_37_G2_G2/B_notx[0] ), .out(\mat_mul/mult_37_G2_G2/ab[1][0] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN2_0_7  ( .a(\mat_mul/mult_37_G2_G2/A_notx[0] ), 
        .b(\mat_mul/mult_37_G2_G2/B_not [7]), .out(
        \mat_mul/mult_37_G2_G2/ab[0][7] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_0_6  ( .a(\mat_mul/mult_37_G2_G2/A_notx[0] ), 
        .b(\mat_mul/mult_37_G2_G2/B_not [6]), .out(
        \mat_mul/mult_37_G2_G2/ab[0][6] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_0_5  ( .a(\mat_mul/mult_37_G2_G2/A_notx[0] ), 
        .b(\mat_mul/mult_37_G2_G2/B_not [5]), .out(
        \mat_mul/mult_37_G2_G2/ab[0][5] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_0_4  ( .a(\mat_mul/mult_37_G2_G2/A_notx[0] ), 
        .b(\mat_mul/mult_37_G2_G2/B_not [4]), .out(
        \mat_mul/mult_37_G2_G2/ab[0][4] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_0_3  ( .a(\mat_mul/mult_37_G2_G2/A_notx[0] ), 
        .b(\mat_mul/mult_37_G2_G2/B_not [3]), .out(
        \mat_mul/mult_37_G2_G2/ab[0][3] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_0_2  ( .a(\mat_mul/mult_37_G2_G2/A_notx[0] ), 
        .b(\mat_mul/mult_37_G2_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2/ab[0][2] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_0_1  ( .a(\mat_mul/mult_37_G2_G2/A_notx[0] ), 
        .b(\mat_mul/mult_37_G2_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2/ab[0][1] ) );
  nor2 \mat_mul/mult_37_G2_G2/AN1_0_0_0  ( .a(
        \mat_mul/mult_37_G2_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G2/B_notx[0] ), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[0] ) );
  inv \mat_mul/mult_37_G2_G2_G2/AN1_7  ( .in(A[7]), .out(
        \mat_mul/mult_37_G2_G2_G2/A_not [7]) );
  inv \mat_mul/mult_37_G2_G2_G2/AN1_6  ( .in(A[6]), .out(
        \mat_mul/mult_37_G2_G2_G2/A_not [6]) );
  inv \mat_mul/mult_37_G2_G2_G2/AN1_5  ( .in(A[5]), .out(
        \mat_mul/mult_37_G2_G2_G2/A_not [5]) );
  inv \mat_mul/mult_37_G2_G2_G2/AN1_4  ( .in(A[4]), .out(
        \mat_mul/mult_37_G2_G2_G2/A_not [4]) );
  inv \mat_mul/mult_37_G2_G2_G2/AN1_3  ( .in(A[3]), .out(
        \mat_mul/mult_37_G2_G2_G2/A_not [3]) );
  inv \mat_mul/mult_37_G2_G2_G2/AN1_2  ( .in(A[2]), .out(
        \mat_mul/mult_37_G2_G2_G2/A_not [2]) );
  inv \mat_mul/mult_37_G2_G2_G2/AN1_1  ( .in(A[1]), .out(
        \mat_mul/mult_37_G2_G2_G2/A_not [1]) );
  inv \mat_mul/mult_37_G2_G2_G2/AN1_0  ( .in(A[0]), .out(
        \mat_mul/mult_37_G2_G2_G2/A_notx[0] ) );
  inv \mat_mul/mult_37_G2_G2_G2/AN1_7_0  ( .in(\mat_add/r106/B_AS [7]), .out(
        \mat_mul/mult_37_G2_G2_G2/B_not [7]) );
  inv \mat_mul/mult_37_G2_G2_G2/AN1_6_0  ( .in(\mat_add/r106/B_AS [6]), .out(
        \mat_mul/mult_37_G2_G2_G2/B_not [6]) );
  inv \mat_mul/mult_37_G2_G2_G2/AN1_5_0  ( .in(\mat_add/r106/B_AS [5]), .out(
        \mat_mul/mult_37_G2_G2_G2/B_not [5]) );
  inv \mat_mul/mult_37_G2_G2_G2/AN1_4_0  ( .in(\mat_add/r106/B_AS [4]), .out(
        \mat_mul/mult_37_G2_G2_G2/B_not [4]) );
  inv \mat_mul/mult_37_G2_G2_G2/AN1_3_0  ( .in(\mat_add/r106/B_AS [3]), .out(
        \mat_mul/mult_37_G2_G2_G2/B_not [3]) );
  inv \mat_mul/mult_37_G2_G2_G2/AN1_2_0  ( .in(\mat_add/r106/B_AS [2]), .out(
        \mat_mul/mult_37_G2_G2_G2/B_not [2]) );
  inv \mat_mul/mult_37_G2_G2_G2/AN1_1_0  ( .in(\mat_add/r106/B_AS [1]), .out(
        \mat_mul/mult_37_G2_G2_G2/B_not [1]) );
  inv \mat_mul/mult_37_G2_G2_G2/AN1_0_0  ( .in(\mat_add/r106/B_AS [0]), .out(
        \mat_mul/mult_37_G2_G2_G2/B_notx[0] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN3_7_0  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [7]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[7][0] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_6_1  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [6]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[6][1] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_6_0_0  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [6]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[6][0] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_5_2  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [5]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[5][2] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_5_1  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [5]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[5][1] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_5_0_0  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [5]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[5][0] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_4_3  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [4]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [3]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[4][3] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_4_2  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [4]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[4][2] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_4_1  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [4]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[4][1] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_4_0_0  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [4]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[4][0] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_3_4  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [3]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [4]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[3][4] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_3_3  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [3]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [3]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[3][3] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_3_2  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [3]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[3][2] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_3_1  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [3]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[3][1] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_3_0_0  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [3]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[3][0] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_2_5  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [5]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[2][5] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_2_4  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [4]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[2][4] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_2_3  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [3]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[2][3] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_2_2  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[2][2] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_2_1  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[2][1] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_2_0_0  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [2]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[2][0] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_1_6  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [6]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[1][6] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_1_5  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [5]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[1][5] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_1_4  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [4]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[1][4] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_1_3  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [3]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[1][3] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_1_2  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[1][2] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_1_1  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[1][1] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_1_0_0  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_not [1]), .b(
        \mat_mul/mult_37_G2_G2_G2/B_notx[0] ), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[1][0] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN2_0_7  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [7]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[0][7] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_0_6  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [6]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[0][6] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_0_5  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [5]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[0][5] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_0_4  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [4]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[0][4] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_0_3  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [3]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[0][3] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_0_2  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [2]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[0][2] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_0_1  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G2_G2/B_not [1]), .out(
        \mat_mul/mult_37_G2_G2_G2/ab[0][1] ) );
  nor2 \mat_mul/mult_37_G2_G2_G2/AN1_0_0_0  ( .a(
        \mat_mul/mult_37_G2_G2_G2/A_notx[0] ), .b(
        \mat_mul/mult_37_G2_G2_G2/B_notx[0] ), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[0] ) );
  inv U293 ( .in(\mat_add/r106/B_AS [7]), .out(\mat_sub/r106/B_AS [7]) );
  inv U294 ( .in(\mat_add/r106/B_AS [6]), .out(\mat_sub/r106/B_AS [6]) );
  inv U295 ( .in(\mat_add/r106/B_AS [5]), .out(\mat_sub/r106/B_AS [5]) );
  inv U296 ( .in(\mat_add/r106/B_AS [4]), .out(\mat_sub/r106/B_AS [4]) );
  inv U297 ( .in(\mat_add/r106/B_AS [3]), .out(\mat_sub/r106/B_AS [3]) );
  inv U298 ( .in(\mat_add/r106/B_AS [2]), .out(\mat_sub/r106/B_AS [2]) );
  inv U299 ( .in(\mat_add/r106/B_AS [1]), .out(\mat_sub/r106/B_AS [1]) );
  inv U300 ( .in(\mat_add/r106/B_AS [0]), .out(\mat_sub/r106/B_AS [0]) );
  inv U301 ( .in(\mat_add/r94/B_AS [7]), .out(\mat_sub/r94/B_AS [7]) );
  inv U302 ( .in(\mat_add/r94/B_AS [6]), .out(\mat_sub/r94/B_AS [6]) );
  inv U303 ( .in(\mat_add/r94/B_AS [5]), .out(\mat_sub/r94/B_AS [5]) );
  inv U304 ( .in(\mat_add/r94/B_AS [4]), .out(\mat_sub/r94/B_AS [4]) );
  inv U305 ( .in(\mat_add/r94/B_AS [3]), .out(\mat_sub/r94/B_AS [3]) );
  inv U306 ( .in(\mat_add/r94/B_AS [2]), .out(\mat_sub/r94/B_AS [2]) );
  inv U307 ( .in(\mat_add/r94/B_AS [1]), .out(\mat_sub/r94/B_AS [1]) );
  inv U308 ( .in(\mat_add/r94/B_AS [0]), .out(\mat_sub/r94/B_AS [0]) );
  inv U309 ( .in(\mat_add/r102/B_AS [7]), .out(\mat_sub/r102/B_AS [7]) );
  inv U310 ( .in(\mat_add/r102/B_AS [6]), .out(\mat_sub/r102/B_AS [6]) );
  inv U311 ( .in(\mat_add/r102/B_AS [5]), .out(\mat_sub/r102/B_AS [5]) );
  inv U312 ( .in(\mat_add/r102/B_AS [4]), .out(\mat_sub/r102/B_AS [4]) );
  inv U313 ( .in(\mat_add/r102/B_AS [3]), .out(\mat_sub/r102/B_AS [3]) );
  inv U314 ( .in(\mat_add/r102/B_AS [2]), .out(\mat_sub/r102/B_AS [2]) );
  inv U315 ( .in(\mat_add/r102/B_AS [1]), .out(\mat_sub/r102/B_AS [1]) );
  inv U316 ( .in(\mat_add/r102/B_AS [0]), .out(\mat_sub/r102/B_AS [0]) );
  inv U317 ( .in(\mat_add/r98/B_AS [7]), .out(\mat_sub/r98/B_AS [7]) );
  inv U318 ( .in(\mat_add/r98/B_AS [6]), .out(\mat_sub/r98/B_AS [6]) );
  inv U319 ( .in(\mat_add/r98/B_AS [5]), .out(\mat_sub/r98/B_AS [5]) );
  inv U320 ( .in(\mat_add/r98/B_AS [4]), .out(\mat_sub/r98/B_AS [4]) );
  inv U321 ( .in(\mat_add/r98/B_AS [3]), .out(\mat_sub/r98/B_AS [3]) );
  inv U322 ( .in(\mat_add/r98/B_AS [2]), .out(\mat_sub/r98/B_AS [2]) );
  inv U323 ( .in(\mat_add/r98/B_AS [1]), .out(\mat_sub/r98/B_AS [1]) );
  inv U324 ( .in(\mat_add/r98/B_AS [0]), .out(\mat_sub/r98/B_AS [0]) );
  inv U325 ( .in(n3126), .out(\mat_mul/mult_37_G2_G2_G2/FS_1/TEMP_P[0][0][0] )
         );
  inv U326 ( .in(n3138), .out(\mat_mul/mult_37_G2_G2/FS_1/TEMP_P[0][0][0] ) );
  inv U327 ( .in(n3150), .out(\mat_mul/mult_37_G2_G1_G2/FS_1/TEMP_P[0][0][0] )
         );
  inv U328 ( .in(n3162), .out(\mat_mul/mult_37_G2/FS_1/TEMP_P[0][0][0] ) );
  inv U329 ( .in(n3174), .out(\mat_mul/mult_37_G2_G2_G1/FS_1/TEMP_P[0][0][0] )
         );
  inv U330 ( .in(n3186), .out(\mat_mul/mult_37_G2_G1/FS_1/TEMP_P[0][0][0] ) );
  inv U331 ( .in(n3198), .out(\mat_mul/mult_37_G2_G1_G1/FS_1/TEMP_P[0][0][0] )
         );
  inv U332 ( .in(n3210), .out(\mat_mul/mult_37/FS_1/TEMP_P[0][0][0] ) );
  inv U333 ( .in(n3222), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/FS_1/TEMP_P[0][0][0] ) );
  inv U334 ( .in(n3234), .out(\mat_kron/mult_40_G2_G2_G2/FS_1/TEMP_P[0][0][0] ) );
  inv U335 ( .in(n3246), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/FS_1/TEMP_P[0][0][0] ) );
  inv U336 ( .in(n3258), .out(\mat_kron/mult_40_G2_G2/FS_1/TEMP_P[0][0][0] )
         );
  inv U337 ( .in(n3270), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/FS_1/TEMP_P[0][0][0] ) );
  inv U338 ( .in(n3282), .out(\mat_kron/mult_40_G2_G1_G2/FS_1/TEMP_P[0][0][0] ) );
  inv U339 ( .in(n3294), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/FS_1/TEMP_P[0][0][0] ) );
  inv U340 ( .in(n3306), .out(\mat_kron/mult_40_G2/FS_1/TEMP_P[0][0][0] ) );
  inv U341 ( .in(n3318), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/FS_1/TEMP_P[0][0][0] ) );
  inv U342 ( .in(n3330), .out(\mat_kron/mult_40_G2_G2_G1/FS_1/TEMP_P[0][0][0] ) );
  inv U343 ( .in(n3342), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/FS_1/TEMP_P[0][0][0] ) );
  inv U344 ( .in(n3354), .out(\mat_kron/mult_40_G2_G1/FS_1/TEMP_P[0][0][0] )
         );
  inv U345 ( .in(n3366), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/FS_1/TEMP_P[0][0][0] ) );
  inv U346 ( .in(n3378), .out(\mat_kron/mult_40_G2_G1_G1/FS_1/TEMP_P[0][0][0] ) );
  inv U347 ( .in(n3390), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/FS_1/TEMP_P[0][0][0] ) );
  inv U348 ( .in(n3402), .out(\mat_kron/mult_40/FS_1/TEMP_P[0][0][0] ) );
  inv U349 ( .in(\mat_kron/mult_40_G2_G2/FS_1/TEMP_P[0][0][0] ), .out(n3259)
         );
  inv U350 ( .in(n3260), .out(\mat_kron/mult_40_G2_G2/FS_1/P[0][0][1] ) );
  inv U351 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/FS_1/TEMP_P[0][0][0] ), .out(
        n3247) );
  inv U352 ( .in(n3248), .out(\mat_kron/mult_40_G2_G1_G2_G2/FS_1/P[0][0][1] )
         );
  inv U353 ( .in(\mat_kron/mult_40_G2_G2_G2/FS_1/TEMP_P[0][0][0] ), .out(n3235) );
  inv U354 ( .in(n3236), .out(\mat_kron/mult_40_G2_G2_G2/FS_1/P[0][0][1] ) );
  inv U355 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/FS_1/TEMP_P[0][0][0] ), .out(
        n3223) );
  inv U356 ( .in(n3224), .out(\mat_kron/mult_40_G2_G2_G2_G2/FS_1/P[0][0][1] )
         );
  inv U357 ( .in(\mat_mul/mult_37_G2_G1_G2/FS_1/TEMP_P[0][0][0] ), .out(n3151)
         );
  inv U358 ( .in(n3152), .out(\mat_mul/mult_37_G2_G1_G2/FS_1/P[0][0][1] ) );
  inv U359 ( .in(\mat_mul/mult_37_G2_G2_G2/FS_1/TEMP_P[0][0][0] ), .out(n3127)
         );
  inv U360 ( .in(n3128), .out(\mat_mul/mult_37_G2_G2_G2/FS_1/P[0][0][1] ) );
  inv U361 ( .in(\mat_kron/mult_40_G2_G2/FS_1/P[0][0][1] ), .out(n3261) );
  inv U362 ( .in(n3262), .out(\mat_kron/mult_40_G2_G2/FS_1/P[0][0][2] ) );
  inv U363 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/FS_1/P[0][0][1] ), .out(n3249)
         );
  inv U364 ( .in(n3250), .out(\mat_kron/mult_40_G2_G1_G2_G2/FS_1/P[0][0][2] )
         );
  inv U365 ( .in(\mat_kron/mult_40_G2_G2_G2/FS_1/P[0][0][1] ), .out(n3237) );
  inv U366 ( .in(n3238), .out(\mat_kron/mult_40_G2_G2_G2/FS_1/P[0][0][2] ) );
  inv U367 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/FS_1/P[0][0][1] ), .out(n3225)
         );
  inv U368 ( .in(n3226), .out(\mat_kron/mult_40_G2_G2_G2_G2/FS_1/P[0][0][2] )
         );
  inv U369 ( .in(\mat_mul/mult_37_G2_G1_G2/FS_1/P[0][0][1] ), .out(n3153) );
  inv U370 ( .in(n3154), .out(\mat_mul/mult_37_G2_G1_G2/FS_1/P[0][0][2] ) );
  inv U371 ( .in(\mat_mul/mult_37_G2_G2_G2/FS_1/P[0][0][1] ), .out(n3129) );
  inv U372 ( .in(n3130), .out(\mat_mul/mult_37_G2_G2_G2/FS_1/P[0][0][2] ) );
  inv U373 ( .in(\mat_kron/mult_40_G2_G2/FS_1/P[0][0][2] ), .out(n3263) );
  inv U374 ( .in(n3264), .out(\mat_kron/mult_40_G2_G2/FS_1/P[0][0][3] ) );
  inv U375 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/FS_1/P[0][0][2] ), .out(n3251)
         );
  inv U376 ( .in(n3252), .out(\mat_kron/mult_40_G2_G1_G2_G2/FS_1/P[0][0][3] )
         );
  inv U377 ( .in(\mat_kron/mult_40_G2_G2_G2/FS_1/P[0][0][2] ), .out(n3239) );
  inv U378 ( .in(n3240), .out(\mat_kron/mult_40_G2_G2_G2/FS_1/P[0][0][3] ) );
  inv U379 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/FS_1/P[0][0][2] ), .out(n3227)
         );
  inv U380 ( .in(n3228), .out(\mat_kron/mult_40_G2_G2_G2_G2/FS_1/P[0][0][3] )
         );
  inv U381 ( .in(\mat_mul/mult_37_G2_G1_G2/FS_1/P[0][0][2] ), .out(n3155) );
  inv U382 ( .in(n3156), .out(\mat_mul/mult_37_G2_G1_G2/FS_1/P[0][0][3] ) );
  inv U383 ( .in(\mat_mul/mult_37_G2_G2_G2/FS_1/P[0][0][2] ), .out(n3131) );
  inv U384 ( .in(n3132), .out(\mat_mul/mult_37_G2_G2_G2/FS_1/P[0][0][3] ) );
  inv U385 ( .in(\mat_kron/mult_40_G2_G2/FS_1/P[0][0][3] ), .out(n3265) );
  inv U386 ( .in(n3266), .out(\mat_kron/mult_40_G2_G2/FS_1/TEMP_P[0][1][0] )
         );
  inv U387 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/FS_1/P[0][0][3] ), .out(n3253)
         );
  inv U388 ( .in(n3254), .out(
        \mat_kron/mult_40_G2_G1_G2_G2/FS_1/TEMP_P[0][1][0] ) );
  inv U389 ( .in(\mat_kron/mult_40_G2_G2_G2/FS_1/P[0][0][3] ), .out(n3241) );
  inv U390 ( .in(n3242), .out(\mat_kron/mult_40_G2_G2_G2/FS_1/TEMP_P[0][1][0] ) );
  inv U391 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/FS_1/P[0][0][3] ), .out(n3229)
         );
  inv U392 ( .in(n3230), .out(
        \mat_kron/mult_40_G2_G2_G2_G2/FS_1/TEMP_P[0][1][0] ) );
  inv U393 ( .in(\mat_mul/mult_37_G2_G1_G2/FS_1/P[0][0][3] ), .out(n3157) );
  inv U394 ( .in(n3158), .out(\mat_mul/mult_37_G2_G1_G2/FS_1/TEMP_P[0][1][0] )
         );
  inv U395 ( .in(\mat_mul/mult_37_G2_G2_G2/FS_1/P[0][0][3] ), .out(n3133) );
  inv U396 ( .in(n3134), .out(\mat_mul/mult_37_G2_G2_G2/FS_1/TEMP_P[0][1][0] )
         );
  inv U397 ( .in(\mat_kron/mult_40_G2_G2/FS_1/TEMP_P[0][1][0] ), .out(n3267)
         );
  inv U398 ( .in(n3268), .out(\mat_kron/mult_40_G2_G2/FS_1/P[0][1][1] ) );
  inv U399 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/FS_1/TEMP_P[0][1][0] ), .out(
        n3255) );
  inv U400 ( .in(n3256), .out(\mat_kron/mult_40_G2_G1_G2_G2/FS_1/P[0][1][1] )
         );
  inv U401 ( .in(\mat_kron/mult_40_G2_G2_G2/FS_1/TEMP_P[0][1][0] ), .out(n3243) );
  inv U402 ( .in(n3244), .out(\mat_kron/mult_40_G2_G2_G2/FS_1/P[0][1][1] ) );
  inv U403 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/FS_1/TEMP_P[0][1][0] ), .out(
        n3231) );
  inv U404 ( .in(n3232), .out(\mat_kron/mult_40_G2_G2_G2_G2/FS_1/P[0][1][1] )
         );
  inv U405 ( .in(\mat_mul/mult_37_G2_G1_G2/FS_1/TEMP_P[0][1][0] ), .out(n3159)
         );
  inv U406 ( .in(n3160), .out(\mat_mul/mult_37_G2_G1_G2/FS_1/P[0][1][1] ) );
  inv U407 ( .in(\mat_mul/mult_37_G2_G2_G2/FS_1/TEMP_P[0][1][0] ), .out(n3135)
         );
  inv U408 ( .in(n3136), .out(\mat_mul/mult_37_G2_G2_G2/FS_1/P[0][1][1] ) );
  inv U409 ( .in(\mat_kron/mult_40_G2_G2/FS_1/P[0][1][1] ), .out(n3269) );
  inv U410 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/FS_1/P[0][1][1] ), .out(n3257)
         );
  inv U411 ( .in(\mat_kron/mult_40_G2_G2_G2/FS_1/P[0][1][1] ), .out(n3245) );
  inv U412 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/FS_1/P[0][1][1] ), .out(n3233)
         );
  inv U413 ( .in(\mat_mul/mult_37_G2_G1_G2/FS_1/P[0][1][1] ), .out(n3161) );
  inv U414 ( .in(\mat_mul/mult_37_G2_G2_G2/FS_1/P[0][1][1] ), .out(n3137) );
  inv U415 ( .in(\mat_kron/mult_40_G2/FS_1/TEMP_P[0][0][0] ), .out(n3307) );
  inv U416 ( .in(n3308), .out(\mat_kron/mult_40_G2/FS_1/P[0][0][1] ) );
  inv U417 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/FS_1/TEMP_P[0][0][0] ), .out(
        n3295) );
  inv U418 ( .in(n3296), .out(\mat_kron/mult_40_G2_G1_G1_G2/FS_1/P[0][0][1] )
         );
  inv U419 ( .in(\mat_kron/mult_40_G2_G1_G2/FS_1/TEMP_P[0][0][0] ), .out(n3283) );
  inv U420 ( .in(n3284), .out(\mat_kron/mult_40_G2_G1_G2/FS_1/P[0][0][1] ) );
  inv U421 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/FS_1/TEMP_P[0][0][0] ), .out(
        n3271) );
  inv U422 ( .in(n3272), .out(\mat_kron/mult_40_G2_G2_G1_G2/FS_1/P[0][0][1] )
         );
  inv U423 ( .in(\mat_mul/mult_37_G2/FS_1/TEMP_P[0][0][0] ), .out(n3163) );
  inv U424 ( .in(n3164), .out(\mat_mul/mult_37_G2/FS_1/P[0][0][1] ) );
  inv U425 ( .in(\mat_mul/mult_37_G2_G2/FS_1/TEMP_P[0][0][0] ), .out(n3139) );
  inv U426 ( .in(n3140), .out(\mat_mul/mult_37_G2_G2/FS_1/P[0][0][1] ) );
  inv U427 ( .in(\mat_kron/mult_40_G2/FS_1/P[0][0][1] ), .out(n3309) );
  inv U428 ( .in(n3310), .out(\mat_kron/mult_40_G2/FS_1/P[0][0][2] ) );
  inv U429 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/FS_1/P[0][0][1] ), .out(n3297)
         );
  inv U430 ( .in(n3298), .out(\mat_kron/mult_40_G2_G1_G1_G2/FS_1/P[0][0][2] )
         );
  inv U431 ( .in(\mat_kron/mult_40_G2_G1_G2/FS_1/P[0][0][1] ), .out(n3285) );
  inv U432 ( .in(n3286), .out(\mat_kron/mult_40_G2_G1_G2/FS_1/P[0][0][2] ) );
  inv U433 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/FS_1/P[0][0][1] ), .out(n3273)
         );
  inv U434 ( .in(n3274), .out(\mat_kron/mult_40_G2_G2_G1_G2/FS_1/P[0][0][2] )
         );
  inv U435 ( .in(\mat_mul/mult_37_G2/FS_1/P[0][0][1] ), .out(n3165) );
  inv U436 ( .in(n3166), .out(\mat_mul/mult_37_G2/FS_1/P[0][0][2] ) );
  inv U437 ( .in(\mat_mul/mult_37_G2_G2/FS_1/P[0][0][1] ), .out(n3141) );
  inv U438 ( .in(n3142), .out(\mat_mul/mult_37_G2_G2/FS_1/P[0][0][2] ) );
  inv U439 ( .in(\mat_kron/mult_40_G2/FS_1/P[0][0][2] ), .out(n3311) );
  inv U440 ( .in(n3312), .out(\mat_kron/mult_40_G2/FS_1/P[0][0][3] ) );
  inv U441 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/FS_1/P[0][0][2] ), .out(n3299)
         );
  inv U442 ( .in(n3300), .out(\mat_kron/mult_40_G2_G1_G1_G2/FS_1/P[0][0][3] )
         );
  inv U443 ( .in(\mat_kron/mult_40_G2_G1_G2/FS_1/P[0][0][2] ), .out(n3287) );
  inv U444 ( .in(n3288), .out(\mat_kron/mult_40_G2_G1_G2/FS_1/P[0][0][3] ) );
  inv U445 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/FS_1/P[0][0][2] ), .out(n3275)
         );
  inv U446 ( .in(n3276), .out(\mat_kron/mult_40_G2_G2_G1_G2/FS_1/P[0][0][3] )
         );
  inv U447 ( .in(\mat_mul/mult_37_G2/FS_1/P[0][0][2] ), .out(n3167) );
  inv U448 ( .in(n3168), .out(\mat_mul/mult_37_G2/FS_1/P[0][0][3] ) );
  inv U449 ( .in(\mat_mul/mult_37_G2_G2/FS_1/P[0][0][2] ), .out(n3143) );
  inv U450 ( .in(n3144), .out(\mat_mul/mult_37_G2_G2/FS_1/P[0][0][3] ) );
  inv U451 ( .in(\mat_kron/mult_40_G2/FS_1/P[0][0][3] ), .out(n3313) );
  inv U452 ( .in(n3314), .out(\mat_kron/mult_40_G2/FS_1/TEMP_P[0][1][0] ) );
  inv U453 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/FS_1/P[0][0][3] ), .out(n3301)
         );
  inv U454 ( .in(n3302), .out(
        \mat_kron/mult_40_G2_G1_G1_G2/FS_1/TEMP_P[0][1][0] ) );
  inv U455 ( .in(\mat_kron/mult_40_G2_G1_G2/FS_1/P[0][0][3] ), .out(n3289) );
  inv U456 ( .in(n3290), .out(\mat_kron/mult_40_G2_G1_G2/FS_1/TEMP_P[0][1][0] ) );
  inv U457 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/FS_1/P[0][0][3] ), .out(n3277)
         );
  inv U458 ( .in(n3278), .out(
        \mat_kron/mult_40_G2_G2_G1_G2/FS_1/TEMP_P[0][1][0] ) );
  inv U459 ( .in(\mat_mul/mult_37_G2/FS_1/P[0][0][3] ), .out(n3169) );
  inv U460 ( .in(n3170), .out(\mat_mul/mult_37_G2/FS_1/TEMP_P[0][1][0] ) );
  inv U461 ( .in(\mat_mul/mult_37_G2_G2/FS_1/P[0][0][3] ), .out(n3145) );
  inv U462 ( .in(n3146), .out(\mat_mul/mult_37_G2_G2/FS_1/TEMP_P[0][1][0] ) );
  inv U463 ( .in(\mat_kron/mult_40_G2/FS_1/TEMP_P[0][1][0] ), .out(n3315) );
  inv U464 ( .in(n3316), .out(\mat_kron/mult_40_G2/FS_1/P[0][1][1] ) );
  inv U465 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/FS_1/TEMP_P[0][1][0] ), .out(
        n3303) );
  inv U466 ( .in(n3304), .out(\mat_kron/mult_40_G2_G1_G1_G2/FS_1/P[0][1][1] )
         );
  inv U467 ( .in(\mat_kron/mult_40_G2_G1_G2/FS_1/TEMP_P[0][1][0] ), .out(n3291) );
  inv U468 ( .in(n3292), .out(\mat_kron/mult_40_G2_G1_G2/FS_1/P[0][1][1] ) );
  inv U469 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/FS_1/TEMP_P[0][1][0] ), .out(
        n3279) );
  inv U470 ( .in(n3280), .out(\mat_kron/mult_40_G2_G2_G1_G2/FS_1/P[0][1][1] )
         );
  inv U471 ( .in(\mat_mul/mult_37_G2/FS_1/TEMP_P[0][1][0] ), .out(n3171) );
  inv U472 ( .in(n3172), .out(\mat_mul/mult_37_G2/FS_1/P[0][1][1] ) );
  inv U473 ( .in(\mat_mul/mult_37_G2_G2/FS_1/TEMP_P[0][1][0] ), .out(n3147) );
  inv U474 ( .in(n3148), .out(\mat_mul/mult_37_G2_G2/FS_1/P[0][1][1] ) );
  inv U475 ( .in(\mat_kron/mult_40_G2/FS_1/P[0][1][1] ), .out(n3317) );
  inv U476 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/FS_1/P[0][1][1] ), .out(n3305)
         );
  inv U477 ( .in(\mat_kron/mult_40_G2_G1_G2/FS_1/P[0][1][1] ), .out(n3293) );
  inv U478 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/FS_1/P[0][1][1] ), .out(n3281)
         );
  inv U479 ( .in(\mat_mul/mult_37_G2/FS_1/P[0][1][1] ), .out(n3173) );
  inv U480 ( .in(\mat_mul/mult_37_G2_G2/FS_1/P[0][1][1] ), .out(n3149) );
  inv U481 ( .in(\mat_kron/mult_40_G2_G1/FS_1/TEMP_P[0][0][0] ), .out(n3355)
         );
  inv U482 ( .in(n3356), .out(\mat_kron/mult_40_G2_G1/FS_1/P[0][0][1] ) );
  inv U483 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/FS_1/TEMP_P[0][0][0] ), .out(
        n3343) );
  inv U484 ( .in(n3344), .out(\mat_kron/mult_40_G2_G1_G2_G1/FS_1/P[0][0][1] )
         );
  inv U485 ( .in(\mat_kron/mult_40_G2_G2_G1/FS_1/TEMP_P[0][0][0] ), .out(n3331) );
  inv U486 ( .in(n3332), .out(\mat_kron/mult_40_G2_G2_G1/FS_1/P[0][0][1] ) );
  inv U487 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/FS_1/TEMP_P[0][0][0] ), .out(
        n3319) );
  inv U488 ( .in(n3320), .out(\mat_kron/mult_40_G2_G2_G2_G1/FS_1/P[0][0][1] )
         );
  inv U489 ( .in(\mat_mul/mult_37_G2_G1_G1/FS_1/TEMP_P[0][0][0] ), .out(n3199)
         );
  inv U490 ( .in(n3200), .out(\mat_mul/mult_37_G2_G1_G1/FS_1/P[0][0][1] ) );
  inv U491 ( .in(\mat_mul/mult_37_G2_G2_G1/FS_1/TEMP_P[0][0][0] ), .out(n3175)
         );
  inv U492 ( .in(n3176), .out(\mat_mul/mult_37_G2_G2_G1/FS_1/P[0][0][1] ) );
  inv U493 ( .in(\mat_kron/mult_40_G2_G1/FS_1/P[0][0][1] ), .out(n3357) );
  inv U494 ( .in(n3358), .out(\mat_kron/mult_40_G2_G1/FS_1/P[0][0][2] ) );
  inv U495 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/FS_1/P[0][0][1] ), .out(n3345)
         );
  inv U496 ( .in(n3346), .out(\mat_kron/mult_40_G2_G1_G2_G1/FS_1/P[0][0][2] )
         );
  inv U497 ( .in(\mat_kron/mult_40_G2_G2_G1/FS_1/P[0][0][1] ), .out(n3333) );
  inv U498 ( .in(n3334), .out(\mat_kron/mult_40_G2_G2_G1/FS_1/P[0][0][2] ) );
  inv U499 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/FS_1/P[0][0][1] ), .out(n3321)
         );
  inv U500 ( .in(n3322), .out(\mat_kron/mult_40_G2_G2_G2_G1/FS_1/P[0][0][2] )
         );
  inv U501 ( .in(\mat_mul/mult_37_G2_G1_G1/FS_1/P[0][0][1] ), .out(n3201) );
  inv U502 ( .in(n3202), .out(\mat_mul/mult_37_G2_G1_G1/FS_1/P[0][0][2] ) );
  inv U503 ( .in(\mat_mul/mult_37_G2_G2_G1/FS_1/P[0][0][1] ), .out(n3177) );
  inv U504 ( .in(n3178), .out(\mat_mul/mult_37_G2_G2_G1/FS_1/P[0][0][2] ) );
  inv U505 ( .in(\mat_kron/mult_40_G2_G1/FS_1/P[0][0][2] ), .out(n3359) );
  inv U506 ( .in(n3360), .out(\mat_kron/mult_40_G2_G1/FS_1/P[0][0][3] ) );
  inv U507 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/FS_1/P[0][0][2] ), .out(n3347)
         );
  inv U508 ( .in(n3348), .out(\mat_kron/mult_40_G2_G1_G2_G1/FS_1/P[0][0][3] )
         );
  inv U509 ( .in(\mat_kron/mult_40_G2_G2_G1/FS_1/P[0][0][2] ), .out(n3335) );
  inv U510 ( .in(n3336), .out(\mat_kron/mult_40_G2_G2_G1/FS_1/P[0][0][3] ) );
  inv U511 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/FS_1/P[0][0][2] ), .out(n3323)
         );
  inv U512 ( .in(n3324), .out(\mat_kron/mult_40_G2_G2_G2_G1/FS_1/P[0][0][3] )
         );
  inv U513 ( .in(\mat_mul/mult_37_G2_G1_G1/FS_1/P[0][0][2] ), .out(n3203) );
  inv U514 ( .in(n3204), .out(\mat_mul/mult_37_G2_G1_G1/FS_1/P[0][0][3] ) );
  inv U515 ( .in(\mat_mul/mult_37_G2_G2_G1/FS_1/P[0][0][2] ), .out(n3179) );
  inv U516 ( .in(n3180), .out(\mat_mul/mult_37_G2_G2_G1/FS_1/P[0][0][3] ) );
  inv U517 ( .in(\mat_kron/mult_40_G2_G1/FS_1/P[0][0][3] ), .out(n3361) );
  inv U518 ( .in(n3362), .out(\mat_kron/mult_40_G2_G1/FS_1/TEMP_P[0][1][0] )
         );
  inv U519 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/FS_1/P[0][0][3] ), .out(n3349)
         );
  inv U520 ( .in(n3350), .out(
        \mat_kron/mult_40_G2_G1_G2_G1/FS_1/TEMP_P[0][1][0] ) );
  inv U521 ( .in(\mat_kron/mult_40_G2_G2_G1/FS_1/P[0][0][3] ), .out(n3337) );
  inv U522 ( .in(n3338), .out(\mat_kron/mult_40_G2_G2_G1/FS_1/TEMP_P[0][1][0] ) );
  inv U523 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/FS_1/P[0][0][3] ), .out(n3325)
         );
  inv U524 ( .in(n3326), .out(
        \mat_kron/mult_40_G2_G2_G2_G1/FS_1/TEMP_P[0][1][0] ) );
  inv U525 ( .in(\mat_mul/mult_37_G2_G1_G1/FS_1/P[0][0][3] ), .out(n3205) );
  inv U526 ( .in(n3206), .out(\mat_mul/mult_37_G2_G1_G1/FS_1/TEMP_P[0][1][0] )
         );
  inv U527 ( .in(\mat_mul/mult_37_G2_G2_G1/FS_1/P[0][0][3] ), .out(n3181) );
  inv U528 ( .in(n3182), .out(\mat_mul/mult_37_G2_G2_G1/FS_1/TEMP_P[0][1][0] )
         );
  inv U529 ( .in(\mat_kron/mult_40_G2_G1/FS_1/TEMP_P[0][1][0] ), .out(n3363)
         );
  inv U530 ( .in(n3364), .out(\mat_kron/mult_40_G2_G1/FS_1/P[0][1][1] ) );
  inv U531 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/FS_1/TEMP_P[0][1][0] ), .out(
        n3351) );
  inv U532 ( .in(n3352), .out(\mat_kron/mult_40_G2_G1_G2_G1/FS_1/P[0][1][1] )
         );
  inv U533 ( .in(\mat_kron/mult_40_G2_G2_G1/FS_1/TEMP_P[0][1][0] ), .out(n3339) );
  inv U534 ( .in(n3340), .out(\mat_kron/mult_40_G2_G2_G1/FS_1/P[0][1][1] ) );
  inv U535 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/FS_1/TEMP_P[0][1][0] ), .out(
        n3327) );
  inv U536 ( .in(n3328), .out(\mat_kron/mult_40_G2_G2_G2_G1/FS_1/P[0][1][1] )
         );
  inv U537 ( .in(\mat_mul/mult_37_G2_G1_G1/FS_1/TEMP_P[0][1][0] ), .out(n3207)
         );
  inv U538 ( .in(n3208), .out(\mat_mul/mult_37_G2_G1_G1/FS_1/P[0][1][1] ) );
  inv U539 ( .in(\mat_mul/mult_37_G2_G2_G1/FS_1/TEMP_P[0][1][0] ), .out(n3183)
         );
  inv U540 ( .in(n3184), .out(\mat_mul/mult_37_G2_G2_G1/FS_1/P[0][1][1] ) );
  inv U541 ( .in(\mat_kron/mult_40_G2_G1/FS_1/P[0][1][1] ), .out(n3365) );
  inv U542 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/FS_1/P[0][1][1] ), .out(n3353)
         );
  inv U543 ( .in(\mat_kron/mult_40_G2_G2_G1/FS_1/P[0][1][1] ), .out(n3341) );
  inv U544 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/FS_1/P[0][1][1] ), .out(n3329)
         );
  inv U545 ( .in(\mat_mul/mult_37_G2_G1_G1/FS_1/P[0][1][1] ), .out(n3209) );
  inv U546 ( .in(\mat_mul/mult_37_G2_G2_G1/FS_1/P[0][1][1] ), .out(n3185) );
  inv U547 ( .in(\mat_kron/mult_40/FS_1/TEMP_P[0][0][0] ), .out(n3403) );
  inv U548 ( .in(n3404), .out(\mat_kron/mult_40/FS_1/P[0][0][1] ) );
  inv U549 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/FS_1/TEMP_P[0][0][0] ), .out(
        n3391) );
  inv U550 ( .in(n3392), .out(\mat_kron/mult_40_G2_G1_G1_G1/FS_1/P[0][0][1] )
         );
  inv U551 ( .in(\mat_kron/mult_40_G2_G1_G1/FS_1/TEMP_P[0][0][0] ), .out(n3379) );
  inv U552 ( .in(n3380), .out(\mat_kron/mult_40_G2_G1_G1/FS_1/P[0][0][1] ) );
  inv U553 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/FS_1/TEMP_P[0][0][0] ), .out(
        n3367) );
  inv U554 ( .in(n3368), .out(\mat_kron/mult_40_G2_G2_G1_G1/FS_1/P[0][0][1] )
         );
  inv U555 ( .in(\mat_mul/mult_37/FS_1/TEMP_P[0][0][0] ), .out(n3211) );
  inv U556 ( .in(n3212), .out(\mat_mul/mult_37/FS_1/P[0][0][1] ) );
  inv U557 ( .in(\mat_mul/mult_37_G2_G1/FS_1/TEMP_P[0][0][0] ), .out(n3187) );
  inv U558 ( .in(n3188), .out(\mat_mul/mult_37_G2_G1/FS_1/P[0][0][1] ) );
  inv U559 ( .in(\mat_kron/mult_40/FS_1/P[0][0][1] ), .out(n3405) );
  inv U560 ( .in(n3406), .out(\mat_kron/mult_40/FS_1/P[0][0][2] ) );
  inv U561 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/FS_1/P[0][0][1] ), .out(n3393)
         );
  inv U562 ( .in(n3394), .out(\mat_kron/mult_40_G2_G1_G1_G1/FS_1/P[0][0][2] )
         );
  inv U563 ( .in(\mat_kron/mult_40_G2_G1_G1/FS_1/P[0][0][1] ), .out(n3381) );
  inv U564 ( .in(n3382), .out(\mat_kron/mult_40_G2_G1_G1/FS_1/P[0][0][2] ) );
  inv U565 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/FS_1/P[0][0][1] ), .out(n3369)
         );
  inv U566 ( .in(n3370), .out(\mat_kron/mult_40_G2_G2_G1_G1/FS_1/P[0][0][2] )
         );
  inv U567 ( .in(\mat_mul/mult_37/FS_1/P[0][0][1] ), .out(n3213) );
  inv U568 ( .in(n3214), .out(\mat_mul/mult_37/FS_1/P[0][0][2] ) );
  inv U569 ( .in(\mat_mul/mult_37_G2_G1/FS_1/P[0][0][1] ), .out(n3189) );
  inv U570 ( .in(n3190), .out(\mat_mul/mult_37_G2_G1/FS_1/P[0][0][2] ) );
  inv U571 ( .in(\mat_kron/mult_40/FS_1/P[0][0][2] ), .out(n3407) );
  inv U572 ( .in(n3408), .out(\mat_kron/mult_40/FS_1/P[0][0][3] ) );
  inv U573 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/FS_1/P[0][0][2] ), .out(n3395)
         );
  inv U574 ( .in(n3396), .out(\mat_kron/mult_40_G2_G1_G1_G1/FS_1/P[0][0][3] )
         );
  inv U575 ( .in(\mat_kron/mult_40_G2_G1_G1/FS_1/P[0][0][2] ), .out(n3383) );
  inv U576 ( .in(n3384), .out(\mat_kron/mult_40_G2_G1_G1/FS_1/P[0][0][3] ) );
  inv U577 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/FS_1/P[0][0][2] ), .out(n3371)
         );
  inv U578 ( .in(n3372), .out(\mat_kron/mult_40_G2_G2_G1_G1/FS_1/P[0][0][3] )
         );
  inv U579 ( .in(\mat_mul/mult_37/FS_1/P[0][0][2] ), .out(n3215) );
  inv U580 ( .in(n3216), .out(\mat_mul/mult_37/FS_1/P[0][0][3] ) );
  inv U581 ( .in(\mat_mul/mult_37_G2_G1/FS_1/P[0][0][2] ), .out(n3191) );
  inv U582 ( .in(n3192), .out(\mat_mul/mult_37_G2_G1/FS_1/P[0][0][3] ) );
  inv U583 ( .in(\mat_kron/mult_40/FS_1/P[0][0][3] ), .out(n3409) );
  inv U584 ( .in(n3410), .out(\mat_kron/mult_40/FS_1/TEMP_P[0][1][0] ) );
  inv U585 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/FS_1/P[0][0][3] ), .out(n3397)
         );
  inv U586 ( .in(n3398), .out(
        \mat_kron/mult_40_G2_G1_G1_G1/FS_1/TEMP_P[0][1][0] ) );
  inv U587 ( .in(\mat_kron/mult_40_G2_G1_G1/FS_1/P[0][0][3] ), .out(n3385) );
  inv U588 ( .in(n3386), .out(\mat_kron/mult_40_G2_G1_G1/FS_1/TEMP_P[0][1][0] ) );
  inv U589 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/FS_1/P[0][0][3] ), .out(n3373)
         );
  inv U590 ( .in(n3374), .out(
        \mat_kron/mult_40_G2_G2_G1_G1/FS_1/TEMP_P[0][1][0] ) );
  inv U591 ( .in(\mat_mul/mult_37/FS_1/P[0][0][3] ), .out(n3217) );
  inv U592 ( .in(n3218), .out(\mat_mul/mult_37/FS_1/TEMP_P[0][1][0] ) );
  inv U593 ( .in(\mat_mul/mult_37_G2_G1/FS_1/P[0][0][3] ), .out(n3193) );
  inv U594 ( .in(n3194), .out(\mat_mul/mult_37_G2_G1/FS_1/TEMP_P[0][1][0] ) );
  inv U595 ( .in(\mat_kron/mult_40/FS_1/TEMP_P[0][1][0] ), .out(n3411) );
  inv U596 ( .in(n3412), .out(\mat_kron/mult_40/FS_1/P[0][1][1] ) );
  inv U597 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/FS_1/TEMP_P[0][1][0] ), .out(
        n3399) );
  inv U598 ( .in(n3400), .out(\mat_kron/mult_40_G2_G1_G1_G1/FS_1/P[0][1][1] )
         );
  inv U599 ( .in(\mat_kron/mult_40_G2_G1_G1/FS_1/TEMP_P[0][1][0] ), .out(n3387) );
  inv U600 ( .in(n3388), .out(\mat_kron/mult_40_G2_G1_G1/FS_1/P[0][1][1] ) );
  inv U601 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/FS_1/TEMP_P[0][1][0] ), .out(
        n3375) );
  inv U602 ( .in(n3376), .out(\mat_kron/mult_40_G2_G2_G1_G1/FS_1/P[0][1][1] )
         );
  inv U603 ( .in(\mat_mul/mult_37/FS_1/TEMP_P[0][1][0] ), .out(n3219) );
  inv U604 ( .in(n3220), .out(\mat_mul/mult_37/FS_1/P[0][1][1] ) );
  inv U605 ( .in(\mat_mul/mult_37_G2_G1/FS_1/TEMP_P[0][1][0] ), .out(n3195) );
  inv U606 ( .in(n3196), .out(\mat_mul/mult_37_G2_G1/FS_1/P[0][1][1] ) );
  inv U607 ( .in(\mat_kron/mult_40/FS_1/P[0][1][1] ), .out(n3413) );
  inv U608 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/FS_1/P[0][1][1] ), .out(n3401)
         );
  inv U609 ( .in(\mat_kron/mult_40_G2_G1_G1/FS_1/P[0][1][1] ), .out(n3389) );
  inv U610 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/FS_1/P[0][1][1] ), .out(n3377)
         );
  inv U611 ( .in(\mat_mul/mult_37/FS_1/P[0][1][1] ), .out(n3221) );
  inv U612 ( .in(\mat_mul/mult_37_G2_G1/FS_1/P[0][1][1] ), .out(n3197) );
  nand2 U613 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[0][6] ), .b(
        \mat_mul/mult_37_G2_G2_G2/ab[1][5] ), .out(n164) );
  nand2 U614 ( .a(\mat_mul/mult_37_G2_G2/ab[0][6] ), .b(
        \mat_mul/mult_37_G2_G2/ab[1][5] ), .out(n165) );
  nand2 U615 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[0][6] ), .b(
        \mat_mul/mult_37_G2_G1_G2/ab[1][5] ), .out(n166) );
  nand2 U616 ( .a(\mat_mul/mult_37_G2/ab[0][6] ), .b(
        \mat_mul/mult_37_G2/ab[1][5] ), .out(n167) );
  nand2 U617 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[0][6] ), .b(
        \mat_mul/mult_37_G2_G2_G1/ab[1][5] ), .out(n168) );
  nand2 U618 ( .a(\mat_mul/mult_37_G2_G1/ab[0][6] ), .b(
        \mat_mul/mult_37_G2_G1/ab[1][5] ), .out(n169) );
  nand2 U619 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[0][6] ), .b(
        \mat_mul/mult_37_G2_G1_G1/ab[1][5] ), .out(n170) );
  nand2 U620 ( .a(\mat_mul/mult_37/ab[0][6] ), .b(\mat_mul/mult_37/ab[1][5] ), 
        .out(n171) );
  nand2 U621 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[0][6] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[1][5] ), .out(n172) );
  nand2 U622 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[0][6] ), .b(
        \mat_kron/mult_40_G2_G2_G2/ab[1][5] ), .out(n173) );
  nand2 U623 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[0][6] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[1][5] ), .out(n174) );
  nand2 U624 ( .a(\mat_kron/mult_40_G2_G2/ab[0][6] ), .b(
        \mat_kron/mult_40_G2_G2/ab[1][5] ), .out(n175) );
  nand2 U625 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[0][6] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[1][5] ), .out(n176) );
  nand2 U626 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[0][6] ), .b(
        \mat_kron/mult_40_G2_G1_G2/ab[1][5] ), .out(n177) );
  nand2 U627 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[0][6] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[1][5] ), .out(n178) );
  nand2 U628 ( .a(\mat_kron/mult_40_G2/ab[0][6] ), .b(
        \mat_kron/mult_40_G2/ab[1][5] ), .out(n179) );
  nand2 U629 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[0][6] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[1][5] ), .out(n180) );
  nand2 U630 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[0][6] ), .b(
        \mat_kron/mult_40_G2_G2_G1/ab[1][5] ), .out(n181) );
  nand2 U631 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[0][6] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[1][5] ), .out(n182) );
  nand2 U632 ( .a(\mat_kron/mult_40_G2_G1/ab[0][6] ), .b(
        \mat_kron/mult_40_G2_G1/ab[1][5] ), .out(n183) );
  nand2 U633 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[0][6] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[1][5] ), .out(n184) );
  nand2 U634 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[0][6] ), .b(
        \mat_kron/mult_40_G2_G1_G1/ab[1][5] ), .out(n185) );
  nand2 U635 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[0][6] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[1][5] ), .out(n186) );
  nand2 U636 ( .a(\mat_kron/mult_40/ab[0][6] ), .b(\mat_kron/mult_40/ab[1][5] ), .out(n187) );
  aoi12 U637 ( .b(\mat_sub/r98/B_AS [0]), .c(A[16]), .a(n189), .out(n188) );
  aoi12 U638 ( .b(\mat_sub/r102/B_AS [0]), .c(A[8]), .a(n191), .out(n190) );
  aoi12 U639 ( .b(\mat_sub/r94/B_AS [0]), .c(A[24]), .a(n193), .out(n192) );
  aoi12 U640 ( .b(\mat_sub/r106/B_AS [0]), .c(A[0]), .a(n195), .out(n194) );
  aoi22 U641 ( .a(n197), .b(n198), .c(\mat_mul/mult_37_G2_G2_G2/ab[2][4] ), 
        .d(n199), .out(n196) );
  nor2 U642 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[2][3] ), .b(n201), .out(n200) );
  aoi22 U643 ( .a(n203), .b(n204), .c(\mat_mul/mult_37_G2_G2_G2/ab[3][3] ), 
        .d(n205), .out(n202) );
  nor2 U644 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[2][2] ), .b(n207), .out(n206) );
  nand2 U645 ( .a(n209), .b(n210), .out(n208) );
  aoi22 U646 ( .a(n212), .b(n213), .c(\mat_mul/mult_37_G2_G2_G2/ab[4][2] ), 
        .d(n214), .out(n211) );
  nand2 U647 ( .a(n216), .b(n217), .out(n215) );
  nor2 U648 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[3][1] ), .b(n219), .out(n218) );
  nor2 U649 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[4][1] ), .b(n221), .out(n220) );
  nor2 U650 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[5][1] ), .b(n223), .out(n222) );
  nand2 U651 ( .a(n225), .b(n226), .out(n224) );
  nand2 U652 ( .a(n228), .b(n229), .out(n227) );
  nand2 U653 ( .a(n231), .b(n232), .out(n230) );
  nor2 U654 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[5][0] ), .b(n234), .out(n233) );
  oai22 U655 ( .a(n236), .b(n237), .c(n238), .d(n239), .out(n235) );
  aoi22 U656 ( .a(n241), .b(n242), .c(\mat_mul/mult_37_G2_G2_G1/ab[2][4] ), 
        .d(n243), .out(n240) );
  nor2 U657 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[2][3] ), .b(n245), .out(n244) );
  aoi22 U658 ( .a(n247), .b(n248), .c(\mat_mul/mult_37_G2_G2_G1/ab[3][3] ), 
        .d(n249), .out(n246) );
  nor2 U659 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[2][2] ), .b(n251), .out(n250) );
  nand2 U660 ( .a(n253), .b(n254), .out(n252) );
  aoi22 U661 ( .a(n256), .b(n257), .c(\mat_mul/mult_37_G2_G2_G1/ab[4][2] ), 
        .d(n258), .out(n255) );
  nand2 U662 ( .a(n260), .b(n261), .out(n259) );
  nor2 U663 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[3][1] ), .b(n263), .out(n262) );
  nor2 U664 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[4][1] ), .b(n265), .out(n264) );
  nor2 U665 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[5][1] ), .b(n267), .out(n266) );
  nand2 U666 ( .a(n269), .b(n270), .out(n268) );
  nand2 U667 ( .a(n272), .b(n273), .out(n271) );
  nand2 U668 ( .a(n275), .b(n276), .out(n274) );
  nor2 U669 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[5][0] ), .b(n278), .out(n277) );
  oai22 U670 ( .a(n280), .b(n281), .c(n282), .d(n283), .out(n279) );
  aoi22 U671 ( .a(n285), .b(n286), .c(\mat_mul/mult_37_G2_G2/ab[2][4] ), .d(
        n287), .out(n284) );
  nor2 U672 ( .a(\mat_mul/mult_37_G2_G2/ab[2][3] ), .b(n289), .out(n288) );
  aoi22 U673 ( .a(n291), .b(n292), .c(\mat_mul/mult_37_G2_G2/ab[3][3] ), .d(
        n293), .out(n290) );
  nor2 U674 ( .a(\mat_mul/mult_37_G2_G2/ab[2][2] ), .b(n295), .out(n294) );
  nand2 U675 ( .a(n297), .b(n298), .out(n296) );
  aoi22 U676 ( .a(n300), .b(n301), .c(\mat_mul/mult_37_G2_G2/ab[4][2] ), .d(
        n302), .out(n299) );
  nand2 U677 ( .a(n304), .b(n305), .out(n303) );
  nor2 U678 ( .a(\mat_mul/mult_37_G2_G2/ab[3][1] ), .b(n307), .out(n306) );
  nor2 U679 ( .a(\mat_mul/mult_37_G2_G2/ab[4][1] ), .b(n309), .out(n308) );
  nor2 U680 ( .a(\mat_mul/mult_37_G2_G2/ab[5][1] ), .b(n311), .out(n310) );
  nand2 U681 ( .a(n313), .b(n314), .out(n312) );
  nand2 U682 ( .a(n316), .b(n317), .out(n315) );
  nand2 U683 ( .a(n319), .b(n320), .out(n318) );
  nor2 U684 ( .a(\mat_mul/mult_37_G2_G2/ab[5][0] ), .b(n322), .out(n321) );
  oai22 U685 ( .a(n324), .b(n325), .c(n326), .d(n327), .out(n323) );
  aoi22 U686 ( .a(n329), .b(n330), .c(\mat_mul/mult_37_G2_G1_G2/ab[2][4] ), 
        .d(n331), .out(n328) );
  nor2 U687 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[2][3] ), .b(n333), .out(n332) );
  aoi22 U688 ( .a(n335), .b(n336), .c(\mat_mul/mult_37_G2_G1_G2/ab[3][3] ), 
        .d(n337), .out(n334) );
  nor2 U689 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[2][2] ), .b(n339), .out(n338) );
  nand2 U690 ( .a(n341), .b(n342), .out(n340) );
  aoi22 U691 ( .a(n344), .b(n345), .c(\mat_mul/mult_37_G2_G1_G2/ab[4][2] ), 
        .d(n346), .out(n343) );
  nand2 U692 ( .a(n348), .b(n349), .out(n347) );
  nor2 U693 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[3][1] ), .b(n351), .out(n350) );
  nor2 U694 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[4][1] ), .b(n353), .out(n352) );
  nor2 U695 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[5][1] ), .b(n355), .out(n354) );
  nand2 U696 ( .a(n357), .b(n358), .out(n356) );
  nand2 U697 ( .a(n360), .b(n361), .out(n359) );
  nand2 U698 ( .a(n363), .b(n364), .out(n362) );
  nor2 U699 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[5][0] ), .b(n366), .out(n365) );
  oai22 U700 ( .a(n368), .b(n369), .c(n370), .d(n371), .out(n367) );
  aoi22 U701 ( .a(n373), .b(n374), .c(\mat_mul/mult_37_G2_G1_G1/ab[2][4] ), 
        .d(n375), .out(n372) );
  nor2 U702 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[2][3] ), .b(n377), .out(n376) );
  aoi22 U703 ( .a(n379), .b(n380), .c(\mat_mul/mult_37_G2_G1_G1/ab[3][3] ), 
        .d(n381), .out(n378) );
  nor2 U704 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[2][2] ), .b(n383), .out(n382) );
  nand2 U705 ( .a(n385), .b(n386), .out(n384) );
  aoi22 U706 ( .a(n388), .b(n389), .c(\mat_mul/mult_37_G2_G1_G1/ab[4][2] ), 
        .d(n390), .out(n387) );
  nand2 U707 ( .a(n392), .b(n393), .out(n391) );
  nor2 U708 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[3][1] ), .b(n395), .out(n394) );
  nor2 U709 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[4][1] ), .b(n397), .out(n396) );
  nor2 U710 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[5][1] ), .b(n399), .out(n398) );
  nand2 U711 ( .a(n401), .b(n402), .out(n400) );
  nand2 U712 ( .a(n404), .b(n405), .out(n403) );
  nand2 U713 ( .a(n407), .b(n408), .out(n406) );
  nor2 U714 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[5][0] ), .b(n410), .out(n409) );
  oai22 U715 ( .a(n412), .b(n413), .c(n414), .d(n415), .out(n411) );
  aoi22 U716 ( .a(n417), .b(n418), .c(\mat_mul/mult_37_G2_G1/ab[2][4] ), .d(
        n419), .out(n416) );
  nor2 U717 ( .a(\mat_mul/mult_37_G2_G1/ab[2][3] ), .b(n421), .out(n420) );
  aoi22 U718 ( .a(n423), .b(n424), .c(\mat_mul/mult_37_G2_G1/ab[3][3] ), .d(
        n425), .out(n422) );
  nor2 U719 ( .a(\mat_mul/mult_37_G2_G1/ab[2][2] ), .b(n427), .out(n426) );
  nand2 U720 ( .a(n429), .b(n430), .out(n428) );
  aoi22 U721 ( .a(n432), .b(n433), .c(\mat_mul/mult_37_G2_G1/ab[4][2] ), .d(
        n434), .out(n431) );
  nand2 U722 ( .a(n436), .b(n437), .out(n435) );
  nor2 U723 ( .a(\mat_mul/mult_37_G2_G1/ab[3][1] ), .b(n439), .out(n438) );
  nor2 U724 ( .a(\mat_mul/mult_37_G2_G1/ab[4][1] ), .b(n441), .out(n440) );
  nor2 U725 ( .a(\mat_mul/mult_37_G2_G1/ab[5][1] ), .b(n443), .out(n442) );
  nand2 U726 ( .a(n445), .b(n446), .out(n444) );
  nand2 U727 ( .a(n448), .b(n449), .out(n447) );
  nand2 U728 ( .a(n451), .b(n452), .out(n450) );
  nor2 U729 ( .a(\mat_mul/mult_37_G2_G1/ab[5][0] ), .b(n454), .out(n453) );
  oai22 U730 ( .a(n456), .b(n457), .c(n458), .d(n459), .out(n455) );
  aoi22 U731 ( .a(n461), .b(n462), .c(\mat_mul/mult_37_G2/ab[2][4] ), .d(n463), 
        .out(n460) );
  nor2 U732 ( .a(\mat_mul/mult_37_G2/ab[2][3] ), .b(n465), .out(n464) );
  aoi22 U733 ( .a(n467), .b(n468), .c(\mat_mul/mult_37_G2/ab[3][3] ), .d(n469), 
        .out(n466) );
  nor2 U734 ( .a(\mat_mul/mult_37_G2/ab[2][2] ), .b(n471), .out(n470) );
  nand2 U735 ( .a(n473), .b(n474), .out(n472) );
  aoi22 U736 ( .a(n476), .b(n477), .c(\mat_mul/mult_37_G2/ab[4][2] ), .d(n478), 
        .out(n475) );
  nand2 U737 ( .a(n480), .b(n481), .out(n479) );
  nor2 U738 ( .a(\mat_mul/mult_37_G2/ab[3][1] ), .b(n483), .out(n482) );
  nor2 U739 ( .a(\mat_mul/mult_37_G2/ab[4][1] ), .b(n485), .out(n484) );
  nor2 U740 ( .a(\mat_mul/mult_37_G2/ab[5][1] ), .b(n487), .out(n486) );
  nand2 U741 ( .a(n489), .b(n490), .out(n488) );
  nand2 U742 ( .a(n492), .b(n493), .out(n491) );
  nand2 U743 ( .a(n495), .b(n496), .out(n494) );
  nor2 U744 ( .a(\mat_mul/mult_37_G2/ab[5][0] ), .b(n498), .out(n497) );
  oai22 U745 ( .a(n500), .b(n501), .c(n502), .d(n503), .out(n499) );
  aoi22 U746 ( .a(n505), .b(n506), .c(\mat_mul/mult_37/ab[2][4] ), .d(n507), 
        .out(n504) );
  nor2 U747 ( .a(\mat_mul/mult_37/ab[2][3] ), .b(n509), .out(n508) );
  aoi22 U748 ( .a(n511), .b(n512), .c(\mat_mul/mult_37/ab[3][3] ), .d(n513), 
        .out(n510) );
  nor2 U749 ( .a(\mat_mul/mult_37/ab[2][2] ), .b(n515), .out(n514) );
  nand2 U750 ( .a(n517), .b(n518), .out(n516) );
  aoi22 U751 ( .a(n520), .b(n521), .c(\mat_mul/mult_37/ab[4][2] ), .d(n522), 
        .out(n519) );
  nand2 U752 ( .a(n524), .b(n525), .out(n523) );
  nor2 U753 ( .a(\mat_mul/mult_37/ab[3][1] ), .b(n527), .out(n526) );
  nor2 U754 ( .a(\mat_mul/mult_37/ab[4][1] ), .b(n529), .out(n528) );
  nor2 U755 ( .a(\mat_mul/mult_37/ab[5][1] ), .b(n531), .out(n530) );
  nand2 U756 ( .a(n533), .b(n534), .out(n532) );
  nand2 U757 ( .a(n536), .b(n537), .out(n535) );
  nand2 U758 ( .a(n539), .b(n540), .out(n538) );
  nor2 U759 ( .a(\mat_mul/mult_37/ab[5][0] ), .b(n542), .out(n541) );
  oai22 U760 ( .a(n544), .b(n545), .c(n546), .d(n547), .out(n543) );
  aoi22 U761 ( .a(n549), .b(n550), .c(\mat_kron/mult_40_G2_G2_G2_G2/ab[2][4] ), 
        .d(n551), .out(n548) );
  nor2 U762 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[2][3] ), .b(n553), .out(n552) );
  aoi22 U763 ( .a(n555), .b(n556), .c(\mat_kron/mult_40_G2_G2_G2_G2/ab[3][3] ), 
        .d(n557), .out(n554) );
  nor2 U764 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[2][2] ), .b(n559), .out(n558) );
  nand2 U765 ( .a(n561), .b(n562), .out(n560) );
  aoi22 U766 ( .a(n564), .b(n565), .c(\mat_kron/mult_40_G2_G2_G2_G2/ab[4][2] ), 
        .d(n566), .out(n563) );
  nand2 U767 ( .a(n568), .b(n569), .out(n567) );
  nor2 U768 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[3][1] ), .b(n571), .out(n570) );
  nor2 U769 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[4][1] ), .b(n573), .out(n572) );
  nor2 U770 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[5][1] ), .b(n575), .out(n574) );
  nand2 U771 ( .a(n577), .b(n578), .out(n576) );
  nand2 U772 ( .a(n580), .b(n581), .out(n579) );
  nand2 U773 ( .a(n583), .b(n584), .out(n582) );
  nor2 U774 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[5][0] ), .b(n586), .out(n585) );
  oai22 U775 ( .a(n588), .b(n589), .c(n590), .d(n591), .out(n587) );
  aoi22 U776 ( .a(n593), .b(n594), .c(\mat_kron/mult_40_G2_G2_G2_G1/ab[2][4] ), 
        .d(n595), .out(n592) );
  nor2 U777 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[2][3] ), .b(n597), .out(n596) );
  aoi22 U778 ( .a(n599), .b(n600), .c(\mat_kron/mult_40_G2_G2_G2_G1/ab[3][3] ), 
        .d(n601), .out(n598) );
  nor2 U779 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[2][2] ), .b(n603), .out(n602) );
  nand2 U780 ( .a(n605), .b(n606), .out(n604) );
  aoi22 U781 ( .a(n608), .b(n609), .c(\mat_kron/mult_40_G2_G2_G2_G1/ab[4][2] ), 
        .d(n610), .out(n607) );
  nand2 U782 ( .a(n612), .b(n613), .out(n611) );
  nor2 U783 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[3][1] ), .b(n615), .out(n614) );
  nor2 U784 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[4][1] ), .b(n617), .out(n616) );
  nor2 U785 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[5][1] ), .b(n619), .out(n618) );
  nand2 U786 ( .a(n621), .b(n622), .out(n620) );
  nand2 U787 ( .a(n624), .b(n625), .out(n623) );
  nand2 U788 ( .a(n627), .b(n628), .out(n626) );
  nor2 U789 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[5][0] ), .b(n630), .out(n629) );
  oai22 U790 ( .a(n632), .b(n633), .c(n634), .d(n635), .out(n631) );
  aoi22 U791 ( .a(n637), .b(n638), .c(\mat_kron/mult_40_G2_G2_G2/ab[2][4] ), 
        .d(n639), .out(n636) );
  nor2 U792 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[2][3] ), .b(n641), .out(n640)
         );
  aoi22 U793 ( .a(n643), .b(n644), .c(\mat_kron/mult_40_G2_G2_G2/ab[3][3] ), 
        .d(n645), .out(n642) );
  nor2 U794 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[2][2] ), .b(n647), .out(n646)
         );
  nand2 U795 ( .a(n649), .b(n650), .out(n648) );
  aoi22 U796 ( .a(n652), .b(n653), .c(\mat_kron/mult_40_G2_G2_G2/ab[4][2] ), 
        .d(n654), .out(n651) );
  nand2 U797 ( .a(n656), .b(n657), .out(n655) );
  nor2 U798 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[3][1] ), .b(n659), .out(n658)
         );
  nor2 U799 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[4][1] ), .b(n661), .out(n660)
         );
  nor2 U800 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[5][1] ), .b(n663), .out(n662)
         );
  nand2 U801 ( .a(n665), .b(n666), .out(n664) );
  nand2 U802 ( .a(n668), .b(n669), .out(n667) );
  nand2 U803 ( .a(n671), .b(n672), .out(n670) );
  nor2 U804 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[5][0] ), .b(n674), .out(n673)
         );
  oai22 U805 ( .a(n676), .b(n677), .c(n678), .d(n679), .out(n675) );
  aoi22 U806 ( .a(n681), .b(n682), .c(\mat_kron/mult_40_G2_G2_G1_G2/ab[2][4] ), 
        .d(n683), .out(n680) );
  nor2 U807 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[2][3] ), .b(n685), .out(n684) );
  aoi22 U808 ( .a(n687), .b(n688), .c(\mat_kron/mult_40_G2_G2_G1_G2/ab[3][3] ), 
        .d(n689), .out(n686) );
  nor2 U809 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[2][2] ), .b(n691), .out(n690) );
  nand2 U810 ( .a(n693), .b(n694), .out(n692) );
  aoi22 U811 ( .a(n696), .b(n697), .c(\mat_kron/mult_40_G2_G2_G1_G2/ab[4][2] ), 
        .d(n698), .out(n695) );
  nand2 U812 ( .a(n700), .b(n701), .out(n699) );
  nor2 U813 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[3][1] ), .b(n703), .out(n702) );
  nor2 U814 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[4][1] ), .b(n705), .out(n704) );
  nor2 U815 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[5][1] ), .b(n707), .out(n706) );
  nand2 U816 ( .a(n709), .b(n710), .out(n708) );
  nand2 U817 ( .a(n712), .b(n713), .out(n711) );
  nand2 U818 ( .a(n715), .b(n716), .out(n714) );
  nor2 U819 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[5][0] ), .b(n718), .out(n717) );
  oai22 U820 ( .a(n720), .b(n721), .c(n722), .d(n723), .out(n719) );
  aoi22 U821 ( .a(n725), .b(n726), .c(\mat_kron/mult_40_G2_G2_G1_G1/ab[2][4] ), 
        .d(n727), .out(n724) );
  nor2 U822 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[2][3] ), .b(n729), .out(n728) );
  aoi22 U823 ( .a(n731), .b(n732), .c(\mat_kron/mult_40_G2_G2_G1_G1/ab[3][3] ), 
        .d(n733), .out(n730) );
  nor2 U824 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[2][2] ), .b(n735), .out(n734) );
  nand2 U825 ( .a(n737), .b(n738), .out(n736) );
  aoi22 U826 ( .a(n740), .b(n741), .c(\mat_kron/mult_40_G2_G2_G1_G1/ab[4][2] ), 
        .d(n742), .out(n739) );
  nand2 U827 ( .a(n744), .b(n745), .out(n743) );
  nor2 U828 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[3][1] ), .b(n747), .out(n746) );
  nor2 U829 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[4][1] ), .b(n749), .out(n748) );
  nor2 U830 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[5][1] ), .b(n751), .out(n750) );
  nand2 U831 ( .a(n753), .b(n754), .out(n752) );
  nand2 U832 ( .a(n756), .b(n757), .out(n755) );
  nand2 U833 ( .a(n759), .b(n760), .out(n758) );
  nor2 U834 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[5][0] ), .b(n762), .out(n761) );
  oai22 U835 ( .a(n764), .b(n765), .c(n766), .d(n767), .out(n763) );
  aoi22 U836 ( .a(n769), .b(n770), .c(\mat_kron/mult_40_G2_G2_G1/ab[2][4] ), 
        .d(n771), .out(n768) );
  nor2 U837 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[2][3] ), .b(n773), .out(n772)
         );
  aoi22 U838 ( .a(n775), .b(n776), .c(\mat_kron/mult_40_G2_G2_G1/ab[3][3] ), 
        .d(n777), .out(n774) );
  nor2 U839 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[2][2] ), .b(n779), .out(n778)
         );
  nand2 U840 ( .a(n781), .b(n782), .out(n780) );
  aoi22 U841 ( .a(n784), .b(n785), .c(\mat_kron/mult_40_G2_G2_G1/ab[4][2] ), 
        .d(n786), .out(n783) );
  nand2 U842 ( .a(n788), .b(n789), .out(n787) );
  nor2 U843 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[3][1] ), .b(n791), .out(n790)
         );
  nor2 U844 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[4][1] ), .b(n793), .out(n792)
         );
  nor2 U845 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[5][1] ), .b(n795), .out(n794)
         );
  nand2 U846 ( .a(n797), .b(n798), .out(n796) );
  nand2 U847 ( .a(n800), .b(n801), .out(n799) );
  nand2 U848 ( .a(n803), .b(n804), .out(n802) );
  nor2 U849 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[5][0] ), .b(n806), .out(n805)
         );
  oai22 U850 ( .a(n808), .b(n809), .c(n810), .d(n811), .out(n807) );
  aoi22 U851 ( .a(n813), .b(n814), .c(\mat_kron/mult_40_G2_G2/ab[2][4] ), .d(
        n815), .out(n812) );
  nor2 U852 ( .a(\mat_kron/mult_40_G2_G2/ab[2][3] ), .b(n817), .out(n816) );
  aoi22 U853 ( .a(n819), .b(n820), .c(\mat_kron/mult_40_G2_G2/ab[3][3] ), .d(
        n821), .out(n818) );
  nor2 U854 ( .a(\mat_kron/mult_40_G2_G2/ab[2][2] ), .b(n823), .out(n822) );
  nand2 U855 ( .a(n825), .b(n826), .out(n824) );
  aoi22 U856 ( .a(n828), .b(n829), .c(\mat_kron/mult_40_G2_G2/ab[4][2] ), .d(
        n830), .out(n827) );
  nand2 U857 ( .a(n832), .b(n833), .out(n831) );
  nor2 U858 ( .a(\mat_kron/mult_40_G2_G2/ab[3][1] ), .b(n835), .out(n834) );
  nor2 U859 ( .a(\mat_kron/mult_40_G2_G2/ab[4][1] ), .b(n837), .out(n836) );
  nor2 U860 ( .a(\mat_kron/mult_40_G2_G2/ab[5][1] ), .b(n839), .out(n838) );
  nand2 U861 ( .a(n841), .b(n842), .out(n840) );
  nand2 U862 ( .a(n844), .b(n845), .out(n843) );
  nand2 U863 ( .a(n847), .b(n848), .out(n846) );
  nor2 U864 ( .a(\mat_kron/mult_40_G2_G2/ab[5][0] ), .b(n850), .out(n849) );
  oai22 U865 ( .a(n852), .b(n853), .c(n854), .d(n855), .out(n851) );
  aoi22 U866 ( .a(n857), .b(n858), .c(\mat_kron/mult_40_G2_G1_G2_G2/ab[2][4] ), 
        .d(n859), .out(n856) );
  nor2 U867 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[2][3] ), .b(n861), .out(n860) );
  aoi22 U868 ( .a(n863), .b(n864), .c(\mat_kron/mult_40_G2_G1_G2_G2/ab[3][3] ), 
        .d(n865), .out(n862) );
  nor2 U869 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[2][2] ), .b(n867), .out(n866) );
  nand2 U870 ( .a(n869), .b(n870), .out(n868) );
  aoi22 U871 ( .a(n872), .b(n873), .c(\mat_kron/mult_40_G2_G1_G2_G2/ab[4][2] ), 
        .d(n874), .out(n871) );
  nand2 U872 ( .a(n876), .b(n877), .out(n875) );
  nor2 U873 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[3][1] ), .b(n879), .out(n878) );
  nor2 U874 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[4][1] ), .b(n881), .out(n880) );
  nor2 U875 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[5][1] ), .b(n883), .out(n882) );
  nand2 U876 ( .a(n885), .b(n886), .out(n884) );
  nand2 U877 ( .a(n888), .b(n889), .out(n887) );
  nand2 U878 ( .a(n891), .b(n892), .out(n890) );
  nor2 U879 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[5][0] ), .b(n894), .out(n893) );
  oai22 U880 ( .a(n896), .b(n897), .c(n898), .d(n899), .out(n895) );
  aoi22 U881 ( .a(n901), .b(n902), .c(\mat_kron/mult_40_G2_G1_G2_G1/ab[2][4] ), 
        .d(n903), .out(n900) );
  nor2 U882 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[2][3] ), .b(n905), .out(n904) );
  aoi22 U883 ( .a(n907), .b(n908), .c(\mat_kron/mult_40_G2_G1_G2_G1/ab[3][3] ), 
        .d(n909), .out(n906) );
  nor2 U884 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[2][2] ), .b(n911), .out(n910) );
  nand2 U885 ( .a(n913), .b(n914), .out(n912) );
  aoi22 U886 ( .a(n916), .b(n917), .c(\mat_kron/mult_40_G2_G1_G2_G1/ab[4][2] ), 
        .d(n918), .out(n915) );
  nand2 U887 ( .a(n920), .b(n921), .out(n919) );
  nor2 U888 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[3][1] ), .b(n923), .out(n922) );
  nor2 U889 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[4][1] ), .b(n925), .out(n924) );
  nor2 U890 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[5][1] ), .b(n927), .out(n926) );
  nand2 U891 ( .a(n929), .b(n930), .out(n928) );
  nand2 U892 ( .a(n932), .b(n933), .out(n931) );
  nand2 U893 ( .a(n935), .b(n936), .out(n934) );
  nor2 U894 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[5][0] ), .b(n938), .out(n937) );
  oai22 U895 ( .a(n940), .b(n941), .c(n942), .d(n943), .out(n939) );
  aoi22 U896 ( .a(n945), .b(n946), .c(\mat_kron/mult_40_G2_G1_G2/ab[2][4] ), 
        .d(n947), .out(n944) );
  nor2 U897 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[2][3] ), .b(n949), .out(n948)
         );
  aoi22 U898 ( .a(n951), .b(n952), .c(\mat_kron/mult_40_G2_G1_G2/ab[3][3] ), 
        .d(n953), .out(n950) );
  nor2 U899 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[2][2] ), .b(n955), .out(n954)
         );
  nand2 U900 ( .a(n957), .b(n958), .out(n956) );
  aoi22 U901 ( .a(n960), .b(n961), .c(\mat_kron/mult_40_G2_G1_G2/ab[4][2] ), 
        .d(n962), .out(n959) );
  nand2 U902 ( .a(n964), .b(n965), .out(n963) );
  nor2 U903 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[3][1] ), .b(n967), .out(n966)
         );
  nor2 U904 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[4][1] ), .b(n969), .out(n968)
         );
  nor2 U905 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[5][1] ), .b(n971), .out(n970)
         );
  nand2 U906 ( .a(n973), .b(n974), .out(n972) );
  nand2 U907 ( .a(n976), .b(n977), .out(n975) );
  nand2 U908 ( .a(n979), .b(n980), .out(n978) );
  nor2 U909 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[5][0] ), .b(n982), .out(n981)
         );
  oai22 U910 ( .a(n984), .b(n985), .c(n986), .d(n987), .out(n983) );
  aoi22 U911 ( .a(n989), .b(n990), .c(\mat_kron/mult_40_G2_G1_G1_G2/ab[2][4] ), 
        .d(n991), .out(n988) );
  nor2 U912 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[2][3] ), .b(n993), .out(n992) );
  aoi22 U913 ( .a(n995), .b(n996), .c(\mat_kron/mult_40_G2_G1_G1_G2/ab[3][3] ), 
        .d(n997), .out(n994) );
  nor2 U914 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[2][2] ), .b(n999), .out(n998) );
  nand2 U915 ( .a(n1001), .b(n1002), .out(n1000) );
  aoi22 U916 ( .a(n1004), .b(n1005), .c(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[4][2] ), .d(n1006), .out(n1003) );
  nand2 U917 ( .a(n1008), .b(n1009), .out(n1007) );
  nor2 U918 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[3][1] ), .b(n1011), .out(
        n1010) );
  nor2 U919 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[4][1] ), .b(n1013), .out(
        n1012) );
  nor2 U920 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[5][1] ), .b(n1015), .out(
        n1014) );
  nand2 U921 ( .a(n1017), .b(n1018), .out(n1016) );
  nand2 U922 ( .a(n1020), .b(n1021), .out(n1019) );
  nand2 U923 ( .a(n1023), .b(n1024), .out(n1022) );
  nor2 U924 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[5][0] ), .b(n1026), .out(
        n1025) );
  oai22 U925 ( .a(n1028), .b(n1029), .c(n1030), .d(n1031), .out(n1027) );
  aoi22 U926 ( .a(n1033), .b(n1034), .c(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[2][4] ), .d(n1035), .out(n1032) );
  nor2 U927 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[2][3] ), .b(n1037), .out(
        n1036) );
  aoi22 U928 ( .a(n1039), .b(n1040), .c(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[3][3] ), .d(n1041), .out(n1038) );
  nor2 U929 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[2][2] ), .b(n1043), .out(
        n1042) );
  nand2 U930 ( .a(n1045), .b(n1046), .out(n1044) );
  aoi22 U931 ( .a(n1048), .b(n1049), .c(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[4][2] ), .d(n1050), .out(n1047) );
  nand2 U932 ( .a(n1052), .b(n1053), .out(n1051) );
  nor2 U933 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[3][1] ), .b(n1055), .out(
        n1054) );
  nor2 U934 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[4][1] ), .b(n1057), .out(
        n1056) );
  nor2 U935 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[5][1] ), .b(n1059), .out(
        n1058) );
  nand2 U936 ( .a(n1061), .b(n1062), .out(n1060) );
  nand2 U937 ( .a(n1064), .b(n1065), .out(n1063) );
  nand2 U938 ( .a(n1067), .b(n1068), .out(n1066) );
  nor2 U939 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[5][0] ), .b(n1070), .out(
        n1069) );
  oai22 U940 ( .a(n1072), .b(n1073), .c(n1074), .d(n1075), .out(n1071) );
  aoi22 U941 ( .a(n1077), .b(n1078), .c(\mat_kron/mult_40_G2_G1_G1/ab[2][4] ), 
        .d(n1079), .out(n1076) );
  nor2 U942 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[2][3] ), .b(n1081), .out(n1080)
         );
  aoi22 U943 ( .a(n1083), .b(n1084), .c(\mat_kron/mult_40_G2_G1_G1/ab[3][3] ), 
        .d(n1085), .out(n1082) );
  nor2 U944 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[2][2] ), .b(n1087), .out(n1086)
         );
  nand2 U945 ( .a(n1089), .b(n1090), .out(n1088) );
  aoi22 U946 ( .a(n1092), .b(n1093), .c(\mat_kron/mult_40_G2_G1_G1/ab[4][2] ), 
        .d(n1094), .out(n1091) );
  nand2 U947 ( .a(n1096), .b(n1097), .out(n1095) );
  nor2 U948 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[3][1] ), .b(n1099), .out(n1098)
         );
  nor2 U949 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[4][1] ), .b(n1101), .out(n1100)
         );
  nor2 U950 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[5][1] ), .b(n1103), .out(n1102)
         );
  nand2 U951 ( .a(n1105), .b(n1106), .out(n1104) );
  nand2 U952 ( .a(n1108), .b(n1109), .out(n1107) );
  nand2 U953 ( .a(n1111), .b(n1112), .out(n1110) );
  nor2 U954 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[5][0] ), .b(n1114), .out(n1113)
         );
  oai22 U955 ( .a(n1116), .b(n1117), .c(n1118), .d(n1119), .out(n1115) );
  aoi22 U956 ( .a(n1121), .b(n1122), .c(\mat_kron/mult_40_G2_G1/ab[2][4] ), 
        .d(n1123), .out(n1120) );
  nor2 U957 ( .a(\mat_kron/mult_40_G2_G1/ab[2][3] ), .b(n1125), .out(n1124) );
  aoi22 U958 ( .a(n1127), .b(n1128), .c(\mat_kron/mult_40_G2_G1/ab[3][3] ), 
        .d(n1129), .out(n1126) );
  nor2 U959 ( .a(\mat_kron/mult_40_G2_G1/ab[2][2] ), .b(n1131), .out(n1130) );
  nand2 U960 ( .a(n1133), .b(n1134), .out(n1132) );
  aoi22 U961 ( .a(n1136), .b(n1137), .c(\mat_kron/mult_40_G2_G1/ab[4][2] ), 
        .d(n1138), .out(n1135) );
  nand2 U962 ( .a(n1140), .b(n1141), .out(n1139) );
  nor2 U963 ( .a(\mat_kron/mult_40_G2_G1/ab[3][1] ), .b(n1143), .out(n1142) );
  nor2 U964 ( .a(\mat_kron/mult_40_G2_G1/ab[4][1] ), .b(n1145), .out(n1144) );
  nor2 U965 ( .a(\mat_kron/mult_40_G2_G1/ab[5][1] ), .b(n1147), .out(n1146) );
  nand2 U966 ( .a(n1149), .b(n1150), .out(n1148) );
  nand2 U967 ( .a(n1152), .b(n1153), .out(n1151) );
  nand2 U968 ( .a(n1155), .b(n1156), .out(n1154) );
  nor2 U969 ( .a(\mat_kron/mult_40_G2_G1/ab[5][0] ), .b(n1158), .out(n1157) );
  oai22 U970 ( .a(n1160), .b(n1161), .c(n1162), .d(n1163), .out(n1159) );
  aoi22 U971 ( .a(n1165), .b(n1166), .c(\mat_kron/mult_40_G2/ab[2][4] ), .d(
        n1167), .out(n1164) );
  nor2 U972 ( .a(\mat_kron/mult_40_G2/ab[2][3] ), .b(n1169), .out(n1168) );
  aoi22 U973 ( .a(n1171), .b(n1172), .c(\mat_kron/mult_40_G2/ab[3][3] ), .d(
        n1173), .out(n1170) );
  nor2 U974 ( .a(\mat_kron/mult_40_G2/ab[2][2] ), .b(n1175), .out(n1174) );
  nand2 U975 ( .a(n1177), .b(n1178), .out(n1176) );
  aoi22 U976 ( .a(n1180), .b(n1181), .c(\mat_kron/mult_40_G2/ab[4][2] ), .d(
        n1182), .out(n1179) );
  nand2 U977 ( .a(n1184), .b(n1185), .out(n1183) );
  nor2 U978 ( .a(\mat_kron/mult_40_G2/ab[3][1] ), .b(n1187), .out(n1186) );
  nor2 U979 ( .a(\mat_kron/mult_40_G2/ab[4][1] ), .b(n1189), .out(n1188) );
  nor2 U980 ( .a(\mat_kron/mult_40_G2/ab[5][1] ), .b(n1191), .out(n1190) );
  nand2 U981 ( .a(n1193), .b(n1194), .out(n1192) );
  nand2 U982 ( .a(n1196), .b(n1197), .out(n1195) );
  nand2 U983 ( .a(n1199), .b(n1200), .out(n1198) );
  nor2 U984 ( .a(\mat_kron/mult_40_G2/ab[5][0] ), .b(n1202), .out(n1201) );
  oai22 U985 ( .a(n1204), .b(n1205), .c(n1206), .d(n1207), .out(n1203) );
  aoi22 U986 ( .a(n1209), .b(n1210), .c(\mat_kron/mult_40/ab[2][4] ), .d(n1211), .out(n1208) );
  nor2 U987 ( .a(\mat_kron/mult_40/ab[2][3] ), .b(n1213), .out(n1212) );
  aoi22 U988 ( .a(n1215), .b(n1216), .c(\mat_kron/mult_40/ab[3][3] ), .d(n1217), .out(n1214) );
  nor2 U989 ( .a(\mat_kron/mult_40/ab[2][2] ), .b(n1219), .out(n1218) );
  nand2 U990 ( .a(n1221), .b(n1222), .out(n1220) );
  aoi22 U991 ( .a(n1224), .b(n1225), .c(\mat_kron/mult_40/ab[4][2] ), .d(n1226), .out(n1223) );
  nand2 U992 ( .a(n1228), .b(n1229), .out(n1227) );
  nor2 U993 ( .a(\mat_kron/mult_40/ab[3][1] ), .b(n1231), .out(n1230) );
  nor2 U994 ( .a(\mat_kron/mult_40/ab[4][1] ), .b(n1233), .out(n1232) );
  nor2 U995 ( .a(\mat_kron/mult_40/ab[5][1] ), .b(n1235), .out(n1234) );
  nand2 U996 ( .a(n1237), .b(n1238), .out(n1236) );
  nand2 U997 ( .a(n1240), .b(n1241), .out(n1239) );
  nand2 U998 ( .a(n1243), .b(n1244), .out(n1242) );
  nor2 U999 ( .a(\mat_kron/mult_40/ab[5][0] ), .b(n1246), .out(n1245) );
  oai22 U1000 ( .a(n1248), .b(n1249), .c(n1250), .d(n1251), .out(n1247) );
  nor2 U1001 ( .a(\mat_sub/r106/B_AS [1]), .b(n1253), .out(n1252) );
  nor2 U1002 ( .a(\mat_sub/r106/B_AS [2]), .b(n1255), .out(n1254) );
  nand2 U1003 ( .a(n1257), .b(n1258), .out(n1256) );
  nor2 U1004 ( .a(\mat_sub/r106/B_AS [4]), .b(n1260), .out(n1259) );
  nand2 U1005 ( .a(n1262), .b(n1263), .out(n1261) );
  aoi22 U1006 ( .a(A[6]), .b(n1265), .c(\mat_sub/r106/B_AS [6]), .d(n1266), 
        .out(n1264) );
  nor2 U1007 ( .a(\mat_sub/r94/B_AS [1]), .b(n1268), .out(n1267) );
  nor2 U1008 ( .a(\mat_sub/r94/B_AS [2]), .b(n1270), .out(n1269) );
  nand2 U1009 ( .a(n1272), .b(n1273), .out(n1271) );
  nor2 U1010 ( .a(\mat_sub/r94/B_AS [4]), .b(n1275), .out(n1274) );
  nand2 U1011 ( .a(n1277), .b(n1278), .out(n1276) );
  aoi22 U1012 ( .a(A[30]), .b(n1280), .c(\mat_sub/r94/B_AS [6]), .d(n1281), 
        .out(n1279) );
  nor2 U1013 ( .a(\mat_sub/r98/B_AS [1]), .b(n1283), .out(n1282) );
  nor2 U1014 ( .a(\mat_sub/r98/B_AS [2]), .b(n1285), .out(n1284) );
  nand2 U1015 ( .a(n1287), .b(n1288), .out(n1286) );
  nor2 U1016 ( .a(\mat_sub/r98/B_AS [4]), .b(n1290), .out(n1289) );
  nand2 U1017 ( .a(n1292), .b(n1293), .out(n1291) );
  aoi22 U1018 ( .a(A[22]), .b(n1295), .c(\mat_sub/r98/B_AS [6]), .d(n1296), 
        .out(n1294) );
  nor2 U1019 ( .a(\mat_sub/r102/B_AS [1]), .b(n1298), .out(n1297) );
  nand2 U1020 ( .a(n1300), .b(n1301), .out(n1299) );
  nand2 U1021 ( .a(n1303), .b(n1304), .out(n1302) );
  nand2 U1022 ( .a(n1306), .b(n1307), .out(n1305) );
  nand2 U1023 ( .a(n1309), .b(n1310), .out(n1308) );
  aoi22 U1024 ( .a(A[14]), .b(n1312), .c(\mat_sub/r102/B_AS [6]), .d(n1313), 
        .out(n1311) );
  nor2 U1025 ( .a(n1315), .b(n1316), .out(n1314) );
  nor2 U1026 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ), .out(n1317) );
  nor2 U1027 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[3] ), .out(n1318) );
  nor2 U1028 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ), .out(n1319) );
  nor2 U1029 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[5] ), .out(n1320) );
  nor2 U1030 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ), .out(n1321) );
  nor2 U1031 ( .a(n1323), .b(n1324), .out(n1322) );
  nor2 U1032 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ), .out(n1325) );
  nor2 U1033 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[3] ), .out(n1326) );
  nor2 U1034 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ), .out(n1327) );
  nor2 U1035 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[5] ), .out(n1328) );
  nor2 U1036 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ), .out(n1329) );
  nor2 U1037 ( .a(n1331), .b(n1332), .out(n1330) );
  nor2 U1038 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ), .out(n1333) );
  nor2 U1039 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[3] ), .out(n1334) );
  nor2 U1040 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ), .out(n1335) );
  nor2 U1041 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[5] ), .out(n1336) );
  nor2 U1042 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ), .out(n1337) );
  nor2 U1043 ( .a(n1339), .b(n1340), .out(n1338) );
  nor2 U1044 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ), .out(n1341) );
  nor2 U1045 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[3] ), .out(n1342) );
  nor2 U1046 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ), .out(n1343) );
  nor2 U1047 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[5] ), .out(n1344) );
  nor2 U1048 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ), .out(n1345) );
  nor2 U1049 ( .a(\mat_add/r106/B_AS [1]), .b(A[1]), .out(n1346) );
  nor2 U1050 ( .a(\mat_add/r106/B_AS [2]), .b(A[2]), .out(n1347) );
  nor2 U1051 ( .a(\mat_add/r106/B_AS [3]), .b(A[3]), .out(n1348) );
  nor2 U1052 ( .a(\mat_add/r106/B_AS [4]), .b(A[4]), .out(n1349) );
  nor2 U1053 ( .a(\mat_add/r106/B_AS [5]), .b(A[5]), .out(n1350) );
  aoi22 U1054 ( .a(n1352), .b(n1353), .c(\mat_add/r106/B_AS [6]), .d(A[6]), 
        .out(n1351) );
  nor2 U1055 ( .a(\mat_add/r94/B_AS [1]), .b(A[25]), .out(n1354) );
  nor2 U1056 ( .a(\mat_add/r94/B_AS [2]), .b(A[26]), .out(n1355) );
  nor2 U1057 ( .a(\mat_add/r94/B_AS [3]), .b(A[27]), .out(n1356) );
  nor2 U1058 ( .a(\mat_add/r94/B_AS [4]), .b(A[28]), .out(n1357) );
  nor2 U1059 ( .a(\mat_add/r94/B_AS [5]), .b(A[29]), .out(n1358) );
  aoi22 U1060 ( .a(n1360), .b(n1361), .c(\mat_add/r94/B_AS [6]), .d(A[30]), 
        .out(n1359) );
  nor2 U1061 ( .a(\mat_add/r98/B_AS [1]), .b(A[17]), .out(n1362) );
  nor2 U1062 ( .a(\mat_add/r98/B_AS [2]), .b(A[18]), .out(n1363) );
  nor2 U1063 ( .a(\mat_add/r98/B_AS [3]), .b(A[19]), .out(n1364) );
  nor2 U1064 ( .a(\mat_add/r98/B_AS [4]), .b(A[20]), .out(n1365) );
  nor2 U1065 ( .a(\mat_add/r98/B_AS [5]), .b(A[21]), .out(n1366) );
  aoi22 U1066 ( .a(n1368), .b(n1369), .c(\mat_add/r98/B_AS [6]), .d(A[22]), 
        .out(n1367) );
  nor2 U1067 ( .a(\mat_add/r102/B_AS [1]), .b(A[9]), .out(n1370) );
  nor2 U1068 ( .a(\mat_add/r102/B_AS [2]), .b(A[10]), .out(n1371) );
  nor2 U1069 ( .a(\mat_add/r102/B_AS [3]), .b(A[11]), .out(n1372) );
  nor2 U1070 ( .a(\mat_add/r102/B_AS [4]), .b(A[12]), .out(n1373) );
  nor2 U1071 ( .a(\mat_add/r102/B_AS [5]), .b(A[13]), .out(n1374) );
  aoi22 U1072 ( .a(n1376), .b(n1377), .c(\mat_add/r102/B_AS [6]), .d(A[14]), 
        .out(n1375) );
  xor2 U1073 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[1][5] ), .b(
        \mat_mul/mult_37_G2_G2_G2/ab[0][6] ), .out(n197) );
  xor2 U1074 ( .a(n1378), .b(n197), .out(n203) );
  xor2 U1075 ( .a(n1380), .b(\mat_mul/mult_37_G2_G2_G2/ab[0][5] ), .out(n1379)
         );
  xor2 U1076 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[1][3] ), .b(
        \mat_mul/mult_37_G2_G2_G2/ab[0][4] ), .out(n1381) );
  xor2 U1077 ( .a(n1383), .b(n1379), .out(n1382) );
  xor2 U1078 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[1][2] ), .b(
        \mat_mul/mult_37_G2_G2_G2/ab[0][3] ), .out(n1384) );
  xor2 U1079 ( .a(n1386), .b(n1381), .out(n1385) );
  xor2 U1080 ( .a(n1388), .b(n212), .out(n1387) );
  xor2 U1081 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[1][1] ), .b(
        \mat_mul/mult_37_G2_G2_G2/ab[0][2] ), .out(n1389) );
  xor2 U1082 ( .a(n1391), .b(n1384), .out(n1390) );
  xor2 U1083 ( .a(n1393), .b(n1394), .out(n1392) );
  xor2 U1084 ( .a(n1395), .b(n1396), .out(\mat_mul/mult_37_G2_G2_G2/A1[5] ) );
  xor2 U1085 ( .a(n1397), .b(n1392), .out(\mat_mul/mult_37_G2_G2_G2/A1[3] ) );
  xor2 U1086 ( .a(n1398), .b(n1390), .out(\mat_mul/mult_37_G2_G2_G2/A1[1] ) );
  xor2 U1087 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[1][5] ), .b(
        \mat_mul/mult_37_G2_G2_G1/ab[0][6] ), .out(n241) );
  xor2 U1088 ( .a(n1399), .b(n241), .out(n247) );
  xor2 U1089 ( .a(n1401), .b(\mat_mul/mult_37_G2_G2_G1/ab[0][5] ), .out(n1400)
         );
  xor2 U1090 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[1][3] ), .b(
        \mat_mul/mult_37_G2_G2_G1/ab[0][4] ), .out(n1402) );
  xor2 U1091 ( .a(n1404), .b(n1400), .out(n1403) );
  xor2 U1092 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[1][2] ), .b(
        \mat_mul/mult_37_G2_G2_G1/ab[0][3] ), .out(n1405) );
  xor2 U1093 ( .a(n1407), .b(n1402), .out(n1406) );
  xor2 U1094 ( .a(n1409), .b(n256), .out(n1408) );
  xor2 U1095 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[1][1] ), .b(
        \mat_mul/mult_37_G2_G2_G1/ab[0][2] ), .out(n1410) );
  xor2 U1096 ( .a(n1412), .b(n1405), .out(n1411) );
  xor2 U1097 ( .a(n1414), .b(n1415), .out(n1413) );
  xor2 U1098 ( .a(n1416), .b(n1417), .out(\mat_mul/mult_37_G2_G2_G1/A1[5] ) );
  xor2 U1099 ( .a(n1418), .b(n1413), .out(\mat_mul/mult_37_G2_G2_G1/A1[3] ) );
  xor2 U1100 ( .a(n1419), .b(n1411), .out(\mat_mul/mult_37_G2_G2_G1/A1[1] ) );
  xor2 U1101 ( .a(\mat_mul/mult_37_G2_G2/ab[1][5] ), .b(
        \mat_mul/mult_37_G2_G2/ab[0][6] ), .out(n285) );
  xor2 U1102 ( .a(n1420), .b(n285), .out(n291) );
  xor2 U1103 ( .a(n1422), .b(\mat_mul/mult_37_G2_G2/ab[0][5] ), .out(n1421) );
  xor2 U1104 ( .a(\mat_mul/mult_37_G2_G2/ab[1][3] ), .b(
        \mat_mul/mult_37_G2_G2/ab[0][4] ), .out(n1423) );
  xor2 U1105 ( .a(n1425), .b(n1421), .out(n1424) );
  xor2 U1106 ( .a(\mat_mul/mult_37_G2_G2/ab[1][2] ), .b(
        \mat_mul/mult_37_G2_G2/ab[0][3] ), .out(n1426) );
  xor2 U1107 ( .a(n1428), .b(n1423), .out(n1427) );
  xor2 U1108 ( .a(n1430), .b(n300), .out(n1429) );
  xor2 U1109 ( .a(\mat_mul/mult_37_G2_G2/ab[1][1] ), .b(
        \mat_mul/mult_37_G2_G2/ab[0][2] ), .out(n1431) );
  xor2 U1110 ( .a(n1433), .b(n1426), .out(n1432) );
  xor2 U1111 ( .a(n1435), .b(n1436), .out(n1434) );
  xor2 U1112 ( .a(n1437), .b(n1438), .out(\mat_mul/mult_37_G2_G2/A1[5] ) );
  xor2 U1113 ( .a(n1439), .b(n1434), .out(\mat_mul/mult_37_G2_G2/A1[3] ) );
  xor2 U1114 ( .a(n1440), .b(n1432), .out(\mat_mul/mult_37_G2_G2/A1[1] ) );
  xor2 U1115 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[1][5] ), .b(
        \mat_mul/mult_37_G2_G1_G2/ab[0][6] ), .out(n329) );
  xor2 U1116 ( .a(n1441), .b(n329), .out(n335) );
  xor2 U1117 ( .a(n1443), .b(\mat_mul/mult_37_G2_G1_G2/ab[0][5] ), .out(n1442)
         );
  xor2 U1118 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[1][3] ), .b(
        \mat_mul/mult_37_G2_G1_G2/ab[0][4] ), .out(n1444) );
  xor2 U1119 ( .a(n1446), .b(n1442), .out(n1445) );
  xor2 U1120 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[1][2] ), .b(
        \mat_mul/mult_37_G2_G1_G2/ab[0][3] ), .out(n1447) );
  xor2 U1121 ( .a(n1449), .b(n1444), .out(n1448) );
  xor2 U1122 ( .a(n1451), .b(n344), .out(n1450) );
  xor2 U1123 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[1][1] ), .b(
        \mat_mul/mult_37_G2_G1_G2/ab[0][2] ), .out(n1452) );
  xor2 U1124 ( .a(n1454), .b(n1447), .out(n1453) );
  xor2 U1125 ( .a(n1456), .b(n1457), .out(n1455) );
  xor2 U1126 ( .a(n1458), .b(n1459), .out(\mat_mul/mult_37_G2_G1_G2/A1[5] ) );
  xor2 U1127 ( .a(n1460), .b(n1455), .out(\mat_mul/mult_37_G2_G1_G2/A1[3] ) );
  xor2 U1128 ( .a(n1461), .b(n1453), .out(\mat_mul/mult_37_G2_G1_G2/A1[1] ) );
  xor2 U1129 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[1][5] ), .b(
        \mat_mul/mult_37_G2_G1_G1/ab[0][6] ), .out(n373) );
  xor2 U1130 ( .a(n1462), .b(n373), .out(n379) );
  xor2 U1131 ( .a(n1464), .b(\mat_mul/mult_37_G2_G1_G1/ab[0][5] ), .out(n1463)
         );
  xor2 U1132 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[1][3] ), .b(
        \mat_mul/mult_37_G2_G1_G1/ab[0][4] ), .out(n1465) );
  xor2 U1133 ( .a(n1467), .b(n1463), .out(n1466) );
  xor2 U1134 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[1][2] ), .b(
        \mat_mul/mult_37_G2_G1_G1/ab[0][3] ), .out(n1468) );
  xor2 U1135 ( .a(n1470), .b(n1465), .out(n1469) );
  xor2 U1136 ( .a(n1472), .b(n388), .out(n1471) );
  xor2 U1137 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[1][1] ), .b(
        \mat_mul/mult_37_G2_G1_G1/ab[0][2] ), .out(n1473) );
  xor2 U1138 ( .a(n1475), .b(n1468), .out(n1474) );
  xor2 U1139 ( .a(n1477), .b(n1478), .out(n1476) );
  xor2 U1140 ( .a(n1479), .b(n1480), .out(\mat_mul/mult_37_G2_G1_G1/A1[5] ) );
  xor2 U1141 ( .a(n1481), .b(n1476), .out(\mat_mul/mult_37_G2_G1_G1/A1[3] ) );
  xor2 U1142 ( .a(n1482), .b(n1474), .out(\mat_mul/mult_37_G2_G1_G1/A1[1] ) );
  xor2 U1143 ( .a(\mat_mul/mult_37_G2_G1/ab[1][5] ), .b(
        \mat_mul/mult_37_G2_G1/ab[0][6] ), .out(n417) );
  xor2 U1144 ( .a(n1483), .b(n417), .out(n423) );
  xor2 U1145 ( .a(n1485), .b(\mat_mul/mult_37_G2_G1/ab[0][5] ), .out(n1484) );
  xor2 U1146 ( .a(\mat_mul/mult_37_G2_G1/ab[1][3] ), .b(
        \mat_mul/mult_37_G2_G1/ab[0][4] ), .out(n1486) );
  xor2 U1147 ( .a(n1488), .b(n1484), .out(n1487) );
  xor2 U1148 ( .a(\mat_mul/mult_37_G2_G1/ab[1][2] ), .b(
        \mat_mul/mult_37_G2_G1/ab[0][3] ), .out(n1489) );
  xor2 U1149 ( .a(n1491), .b(n1486), .out(n1490) );
  xor2 U1150 ( .a(n1493), .b(n432), .out(n1492) );
  xor2 U1151 ( .a(\mat_mul/mult_37_G2_G1/ab[1][1] ), .b(
        \mat_mul/mult_37_G2_G1/ab[0][2] ), .out(n1494) );
  xor2 U1152 ( .a(n1496), .b(n1489), .out(n1495) );
  xor2 U1153 ( .a(n1498), .b(n1499), .out(n1497) );
  xor2 U1154 ( .a(n1500), .b(n1501), .out(\mat_mul/mult_37_G2_G1/A1[5] ) );
  xor2 U1155 ( .a(n1502), .b(n1497), .out(\mat_mul/mult_37_G2_G1/A1[3] ) );
  xor2 U1156 ( .a(n1503), .b(n1495), .out(\mat_mul/mult_37_G2_G1/A1[1] ) );
  xor2 U1157 ( .a(\mat_mul/mult_37_G2/ab[1][5] ), .b(
        \mat_mul/mult_37_G2/ab[0][6] ), .out(n461) );
  xor2 U1158 ( .a(n1504), .b(n461), .out(n467) );
  xor2 U1159 ( .a(n1506), .b(\mat_mul/mult_37_G2/ab[0][5] ), .out(n1505) );
  xor2 U1160 ( .a(\mat_mul/mult_37_G2/ab[1][3] ), .b(
        \mat_mul/mult_37_G2/ab[0][4] ), .out(n1507) );
  xor2 U1161 ( .a(n1509), .b(n1505), .out(n1508) );
  xor2 U1162 ( .a(\mat_mul/mult_37_G2/ab[1][2] ), .b(
        \mat_mul/mult_37_G2/ab[0][3] ), .out(n1510) );
  xor2 U1163 ( .a(n1512), .b(n1507), .out(n1511) );
  xor2 U1164 ( .a(n1514), .b(n476), .out(n1513) );
  xor2 U1165 ( .a(\mat_mul/mult_37_G2/ab[1][1] ), .b(
        \mat_mul/mult_37_G2/ab[0][2] ), .out(n1515) );
  xor2 U1166 ( .a(n1517), .b(n1510), .out(n1516) );
  xor2 U1167 ( .a(n1519), .b(n1520), .out(n1518) );
  xor2 U1168 ( .a(n1521), .b(n1522), .out(\mat_mul/mult_37_G2/A1[5] ) );
  xor2 U1169 ( .a(n1523), .b(n1518), .out(\mat_mul/mult_37_G2/A1[3] ) );
  xor2 U1170 ( .a(n1524), .b(n1516), .out(\mat_mul/mult_37_G2/A1[1] ) );
  xor2 U1171 ( .a(\mat_mul/mult_37/ab[1][5] ), .b(\mat_mul/mult_37/ab[0][6] ), 
        .out(n505) );
  xor2 U1172 ( .a(n1525), .b(n505), .out(n511) );
  xor2 U1173 ( .a(n1527), .b(\mat_mul/mult_37/ab[0][5] ), .out(n1526) );
  xor2 U1174 ( .a(\mat_mul/mult_37/ab[1][3] ), .b(\mat_mul/mult_37/ab[0][4] ), 
        .out(n1528) );
  xor2 U1175 ( .a(n1530), .b(n1526), .out(n1529) );
  xor2 U1176 ( .a(\mat_mul/mult_37/ab[1][2] ), .b(\mat_mul/mult_37/ab[0][3] ), 
        .out(n1531) );
  xor2 U1177 ( .a(n1533), .b(n1528), .out(n1532) );
  xor2 U1178 ( .a(n1535), .b(n520), .out(n1534) );
  xor2 U1179 ( .a(\mat_mul/mult_37/ab[1][1] ), .b(\mat_mul/mult_37/ab[0][2] ), 
        .out(n1536) );
  xor2 U1180 ( .a(n1538), .b(n1531), .out(n1537) );
  xor2 U1181 ( .a(n1540), .b(n1541), .out(n1539) );
  xor2 U1182 ( .a(n1542), .b(n1543), .out(\mat_mul/mult_37/A1[5] ) );
  xor2 U1183 ( .a(n1544), .b(n1539), .out(\mat_mul/mult_37/A1[3] ) );
  xor2 U1184 ( .a(n1545), .b(n1537), .out(\mat_mul/mult_37/A1[1] ) );
  xor2 U1185 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[1][5] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[0][6] ), .out(n549) );
  xor2 U1186 ( .a(n1546), .b(n549), .out(n555) );
  xor2 U1187 ( .a(n1548), .b(\mat_kron/mult_40_G2_G2_G2_G2/ab[0][5] ), .out(
        n1547) );
  xor2 U1188 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[0][4] ), .out(n1549) );
  xor2 U1189 ( .a(n1551), .b(n1547), .out(n1550) );
  xor2 U1190 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[1][2] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[0][3] ), .out(n1552) );
  xor2 U1191 ( .a(n1554), .b(n1549), .out(n1553) );
  xor2 U1192 ( .a(n1556), .b(n564), .out(n1555) );
  xor2 U1193 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[1][1] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[0][2] ), .out(n1557) );
  xor2 U1194 ( .a(n1559), .b(n1552), .out(n1558) );
  xor2 U1195 ( .a(n1561), .b(n1562), .out(n1560) );
  xor2 U1196 ( .a(n1563), .b(n1564), .out(\mat_kron/mult_40_G2_G2_G2_G2/A1[5] ) );
  xor2 U1197 ( .a(n1565), .b(n1560), .out(\mat_kron/mult_40_G2_G2_G2_G2/A1[3] ) );
  xor2 U1198 ( .a(n1566), .b(n1558), .out(\mat_kron/mult_40_G2_G2_G2_G2/A1[1] ) );
  xor2 U1199 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[1][5] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[0][6] ), .out(n593) );
  xor2 U1200 ( .a(n1567), .b(n593), .out(n599) );
  xor2 U1201 ( .a(n1569), .b(\mat_kron/mult_40_G2_G2_G2_G1/ab[0][5] ), .out(
        n1568) );
  xor2 U1202 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[0][4] ), .out(n1570) );
  xor2 U1203 ( .a(n1572), .b(n1568), .out(n1571) );
  xor2 U1204 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[1][2] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[0][3] ), .out(n1573) );
  xor2 U1205 ( .a(n1575), .b(n1570), .out(n1574) );
  xor2 U1206 ( .a(n1577), .b(n608), .out(n1576) );
  xor2 U1207 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[1][1] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[0][2] ), .out(n1578) );
  xor2 U1208 ( .a(n1580), .b(n1573), .out(n1579) );
  xor2 U1209 ( .a(n1582), .b(n1583), .out(n1581) );
  xor2 U1210 ( .a(n1584), .b(n1585), .out(\mat_kron/mult_40_G2_G2_G2_G1/A1[5] ) );
  xor2 U1211 ( .a(n1586), .b(n1581), .out(\mat_kron/mult_40_G2_G2_G2_G1/A1[3] ) );
  xor2 U1212 ( .a(n1587), .b(n1579), .out(\mat_kron/mult_40_G2_G2_G2_G1/A1[1] ) );
  xor2 U1213 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[1][5] ), .b(
        \mat_kron/mult_40_G2_G2_G2/ab[0][6] ), .out(n637) );
  xor2 U1214 ( .a(n1588), .b(n637), .out(n643) );
  xor2 U1215 ( .a(n1590), .b(\mat_kron/mult_40_G2_G2_G2/ab[0][5] ), .out(n1589) );
  xor2 U1216 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G2_G2/ab[0][4] ), .out(n1591) );
  xor2 U1217 ( .a(n1593), .b(n1589), .out(n1592) );
  xor2 U1218 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[1][2] ), .b(
        \mat_kron/mult_40_G2_G2_G2/ab[0][3] ), .out(n1594) );
  xor2 U1219 ( .a(n1596), .b(n1591), .out(n1595) );
  xor2 U1220 ( .a(n1598), .b(n652), .out(n1597) );
  xor2 U1221 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[1][1] ), .b(
        \mat_kron/mult_40_G2_G2_G2/ab[0][2] ), .out(n1599) );
  xor2 U1222 ( .a(n1601), .b(n1594), .out(n1600) );
  xor2 U1223 ( .a(n1603), .b(n1604), .out(n1602) );
  xor2 U1224 ( .a(n1605), .b(n1606), .out(\mat_kron/mult_40_G2_G2_G2/A1[5] )
         );
  xor2 U1225 ( .a(n1607), .b(n1602), .out(\mat_kron/mult_40_G2_G2_G2/A1[3] )
         );
  xor2 U1226 ( .a(n1608), .b(n1600), .out(\mat_kron/mult_40_G2_G2_G2/A1[1] )
         );
  xor2 U1227 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[1][5] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[0][6] ), .out(n681) );
  xor2 U1228 ( .a(n1609), .b(n681), .out(n687) );
  xor2 U1229 ( .a(n1611), .b(\mat_kron/mult_40_G2_G2_G1_G2/ab[0][5] ), .out(
        n1610) );
  xor2 U1230 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[0][4] ), .out(n1612) );
  xor2 U1231 ( .a(n1614), .b(n1610), .out(n1613) );
  xor2 U1232 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[1][2] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[0][3] ), .out(n1615) );
  xor2 U1233 ( .a(n1617), .b(n1612), .out(n1616) );
  xor2 U1234 ( .a(n1619), .b(n696), .out(n1618) );
  xor2 U1235 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[1][1] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[0][2] ), .out(n1620) );
  xor2 U1236 ( .a(n1622), .b(n1615), .out(n1621) );
  xor2 U1237 ( .a(n1624), .b(n1625), .out(n1623) );
  xor2 U1238 ( .a(n1626), .b(n1627), .out(\mat_kron/mult_40_G2_G2_G1_G2/A1[5] ) );
  xor2 U1239 ( .a(n1628), .b(n1623), .out(\mat_kron/mult_40_G2_G2_G1_G2/A1[3] ) );
  xor2 U1240 ( .a(n1629), .b(n1621), .out(\mat_kron/mult_40_G2_G2_G1_G2/A1[1] ) );
  xor2 U1241 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[1][5] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[0][6] ), .out(n725) );
  xor2 U1242 ( .a(n1630), .b(n725), .out(n731) );
  xor2 U1243 ( .a(n1632), .b(\mat_kron/mult_40_G2_G2_G1_G1/ab[0][5] ), .out(
        n1631) );
  xor2 U1244 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[0][4] ), .out(n1633) );
  xor2 U1245 ( .a(n1635), .b(n1631), .out(n1634) );
  xor2 U1246 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[1][2] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[0][3] ), .out(n1636) );
  xor2 U1247 ( .a(n1638), .b(n1633), .out(n1637) );
  xor2 U1248 ( .a(n1640), .b(n740), .out(n1639) );
  xor2 U1249 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[1][1] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[0][2] ), .out(n1641) );
  xor2 U1250 ( .a(n1643), .b(n1636), .out(n1642) );
  xor2 U1251 ( .a(n1645), .b(n1646), .out(n1644) );
  xor2 U1252 ( .a(n1647), .b(n1648), .out(\mat_kron/mult_40_G2_G2_G1_G1/A1[5] ) );
  xor2 U1253 ( .a(n1649), .b(n1644), .out(\mat_kron/mult_40_G2_G2_G1_G1/A1[3] ) );
  xor2 U1254 ( .a(n1650), .b(n1642), .out(\mat_kron/mult_40_G2_G2_G1_G1/A1[1] ) );
  xor2 U1255 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[1][5] ), .b(
        \mat_kron/mult_40_G2_G2_G1/ab[0][6] ), .out(n769) );
  xor2 U1256 ( .a(n1651), .b(n769), .out(n775) );
  xor2 U1257 ( .a(n1653), .b(\mat_kron/mult_40_G2_G2_G1/ab[0][5] ), .out(n1652) );
  xor2 U1258 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G2_G1/ab[0][4] ), .out(n1654) );
  xor2 U1259 ( .a(n1656), .b(n1652), .out(n1655) );
  xor2 U1260 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[1][2] ), .b(
        \mat_kron/mult_40_G2_G2_G1/ab[0][3] ), .out(n1657) );
  xor2 U1261 ( .a(n1659), .b(n1654), .out(n1658) );
  xor2 U1262 ( .a(n1661), .b(n784), .out(n1660) );
  xor2 U1263 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[1][1] ), .b(
        \mat_kron/mult_40_G2_G2_G1/ab[0][2] ), .out(n1662) );
  xor2 U1264 ( .a(n1664), .b(n1657), .out(n1663) );
  xor2 U1265 ( .a(n1666), .b(n1667), .out(n1665) );
  xor2 U1266 ( .a(n1668), .b(n1669), .out(\mat_kron/mult_40_G2_G2_G1/A1[5] )
         );
  xor2 U1267 ( .a(n1670), .b(n1665), .out(\mat_kron/mult_40_G2_G2_G1/A1[3] )
         );
  xor2 U1268 ( .a(n1671), .b(n1663), .out(\mat_kron/mult_40_G2_G2_G1/A1[1] )
         );
  xor2 U1269 ( .a(\mat_kron/mult_40_G2_G2/ab[1][5] ), .b(
        \mat_kron/mult_40_G2_G2/ab[0][6] ), .out(n813) );
  xor2 U1270 ( .a(n1672), .b(n813), .out(n819) );
  xor2 U1271 ( .a(n1674), .b(\mat_kron/mult_40_G2_G2/ab[0][5] ), .out(n1673)
         );
  xor2 U1272 ( .a(\mat_kron/mult_40_G2_G2/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G2/ab[0][4] ), .out(n1675) );
  xor2 U1273 ( .a(n1677), .b(n1673), .out(n1676) );
  xor2 U1274 ( .a(\mat_kron/mult_40_G2_G2/ab[1][2] ), .b(
        \mat_kron/mult_40_G2_G2/ab[0][3] ), .out(n1678) );
  xor2 U1275 ( .a(n1680), .b(n1675), .out(n1679) );
  xor2 U1276 ( .a(n1682), .b(n828), .out(n1681) );
  xor2 U1277 ( .a(\mat_kron/mult_40_G2_G2/ab[1][1] ), .b(
        \mat_kron/mult_40_G2_G2/ab[0][2] ), .out(n1683) );
  xor2 U1278 ( .a(n1685), .b(n1678), .out(n1684) );
  xor2 U1279 ( .a(n1687), .b(n1688), .out(n1686) );
  xor2 U1280 ( .a(n1689), .b(n1690), .out(\mat_kron/mult_40_G2_G2/A1[5] ) );
  xor2 U1281 ( .a(n1691), .b(n1686), .out(\mat_kron/mult_40_G2_G2/A1[3] ) );
  xor2 U1282 ( .a(n1692), .b(n1684), .out(\mat_kron/mult_40_G2_G2/A1[1] ) );
  xor2 U1283 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[1][5] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[0][6] ), .out(n857) );
  xor2 U1284 ( .a(n1693), .b(n857), .out(n863) );
  xor2 U1285 ( .a(n1695), .b(\mat_kron/mult_40_G2_G1_G2_G2/ab[0][5] ), .out(
        n1694) );
  xor2 U1286 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[0][4] ), .out(n1696) );
  xor2 U1287 ( .a(n1698), .b(n1694), .out(n1697) );
  xor2 U1288 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[1][2] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[0][3] ), .out(n1699) );
  xor2 U1289 ( .a(n1701), .b(n1696), .out(n1700) );
  xor2 U1290 ( .a(n1703), .b(n872), .out(n1702) );
  xor2 U1291 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[1][1] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[0][2] ), .out(n1704) );
  xor2 U1292 ( .a(n1706), .b(n1699), .out(n1705) );
  xor2 U1293 ( .a(n1708), .b(n1709), .out(n1707) );
  xor2 U1294 ( .a(n1710), .b(n1711), .out(\mat_kron/mult_40_G2_G1_G2_G2/A1[5] ) );
  xor2 U1295 ( .a(n1712), .b(n1707), .out(\mat_kron/mult_40_G2_G1_G2_G2/A1[3] ) );
  xor2 U1296 ( .a(n1713), .b(n1705), .out(\mat_kron/mult_40_G2_G1_G2_G2/A1[1] ) );
  xor2 U1297 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[1][5] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[0][6] ), .out(n901) );
  xor2 U1298 ( .a(n1714), .b(n901), .out(n907) );
  xor2 U1299 ( .a(n1716), .b(\mat_kron/mult_40_G2_G1_G2_G1/ab[0][5] ), .out(
        n1715) );
  xor2 U1300 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[0][4] ), .out(n1717) );
  xor2 U1301 ( .a(n1719), .b(n1715), .out(n1718) );
  xor2 U1302 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[1][2] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[0][3] ), .out(n1720) );
  xor2 U1303 ( .a(n1722), .b(n1717), .out(n1721) );
  xor2 U1304 ( .a(n1724), .b(n916), .out(n1723) );
  xor2 U1305 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[1][1] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[0][2] ), .out(n1725) );
  xor2 U1306 ( .a(n1727), .b(n1720), .out(n1726) );
  xor2 U1307 ( .a(n1729), .b(n1730), .out(n1728) );
  xor2 U1308 ( .a(n1731), .b(n1732), .out(\mat_kron/mult_40_G2_G1_G2_G1/A1[5] ) );
  xor2 U1309 ( .a(n1733), .b(n1728), .out(\mat_kron/mult_40_G2_G1_G2_G1/A1[3] ) );
  xor2 U1310 ( .a(n1734), .b(n1726), .out(\mat_kron/mult_40_G2_G1_G2_G1/A1[1] ) );
  xor2 U1311 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[1][5] ), .b(
        \mat_kron/mult_40_G2_G1_G2/ab[0][6] ), .out(n945) );
  xor2 U1312 ( .a(n1735), .b(n945), .out(n951) );
  xor2 U1313 ( .a(n1737), .b(\mat_kron/mult_40_G2_G1_G2/ab[0][5] ), .out(n1736) );
  xor2 U1314 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G1_G2/ab[0][4] ), .out(n1738) );
  xor2 U1315 ( .a(n1740), .b(n1736), .out(n1739) );
  xor2 U1316 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[1][2] ), .b(
        \mat_kron/mult_40_G2_G1_G2/ab[0][3] ), .out(n1741) );
  xor2 U1317 ( .a(n1743), .b(n1738), .out(n1742) );
  xor2 U1318 ( .a(n1745), .b(n960), .out(n1744) );
  xor2 U1319 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[1][1] ), .b(
        \mat_kron/mult_40_G2_G1_G2/ab[0][2] ), .out(n1746) );
  xor2 U1320 ( .a(n1748), .b(n1741), .out(n1747) );
  xor2 U1321 ( .a(n1750), .b(n1751), .out(n1749) );
  xor2 U1322 ( .a(n1752), .b(n1753), .out(\mat_kron/mult_40_G2_G1_G2/A1[5] )
         );
  xor2 U1323 ( .a(n1754), .b(n1749), .out(\mat_kron/mult_40_G2_G1_G2/A1[3] )
         );
  xor2 U1324 ( .a(n1755), .b(n1747), .out(\mat_kron/mult_40_G2_G1_G2/A1[1] )
         );
  xor2 U1325 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[1][5] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[0][6] ), .out(n989) );
  xor2 U1326 ( .a(n1756), .b(n989), .out(n995) );
  xor2 U1327 ( .a(n1758), .b(\mat_kron/mult_40_G2_G1_G1_G2/ab[0][5] ), .out(
        n1757) );
  xor2 U1328 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[0][4] ), .out(n1759) );
  xor2 U1329 ( .a(n1761), .b(n1757), .out(n1760) );
  xor2 U1330 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[1][2] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[0][3] ), .out(n1762) );
  xor2 U1331 ( .a(n1764), .b(n1759), .out(n1763) );
  xor2 U1332 ( .a(n1766), .b(n1004), .out(n1765) );
  xor2 U1333 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[1][1] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[0][2] ), .out(n1767) );
  xor2 U1334 ( .a(n1769), .b(n1762), .out(n1768) );
  xor2 U1335 ( .a(n1771), .b(n1772), .out(n1770) );
  xor2 U1336 ( .a(n1773), .b(n1774), .out(\mat_kron/mult_40_G2_G1_G1_G2/A1[5] ) );
  xor2 U1337 ( .a(n1775), .b(n1770), .out(\mat_kron/mult_40_G2_G1_G1_G2/A1[3] ) );
  xor2 U1338 ( .a(n1776), .b(n1768), .out(\mat_kron/mult_40_G2_G1_G1_G2/A1[1] ) );
  xor2 U1339 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[1][5] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[0][6] ), .out(n1033) );
  xor2 U1340 ( .a(n1777), .b(n1033), .out(n1039) );
  xor2 U1341 ( .a(n1779), .b(\mat_kron/mult_40_G2_G1_G1_G1/ab[0][5] ), .out(
        n1778) );
  xor2 U1342 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[0][4] ), .out(n1780) );
  xor2 U1343 ( .a(n1782), .b(n1778), .out(n1781) );
  xor2 U1344 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[1][2] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[0][3] ), .out(n1783) );
  xor2 U1345 ( .a(n1785), .b(n1780), .out(n1784) );
  xor2 U1346 ( .a(n1787), .b(n1048), .out(n1786) );
  xor2 U1347 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[1][1] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[0][2] ), .out(n1788) );
  xor2 U1348 ( .a(n1790), .b(n1783), .out(n1789) );
  xor2 U1349 ( .a(n1792), .b(n1793), .out(n1791) );
  xor2 U1350 ( .a(n1794), .b(n1795), .out(\mat_kron/mult_40_G2_G1_G1_G1/A1[5] ) );
  xor2 U1351 ( .a(n1796), .b(n1791), .out(\mat_kron/mult_40_G2_G1_G1_G1/A1[3] ) );
  xor2 U1352 ( .a(n1797), .b(n1789), .out(\mat_kron/mult_40_G2_G1_G1_G1/A1[1] ) );
  xor2 U1353 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[1][5] ), .b(
        \mat_kron/mult_40_G2_G1_G1/ab[0][6] ), .out(n1077) );
  xor2 U1354 ( .a(n1798), .b(n1077), .out(n1083) );
  xor2 U1355 ( .a(n1800), .b(\mat_kron/mult_40_G2_G1_G1/ab[0][5] ), .out(n1799) );
  xor2 U1356 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G1_G1/ab[0][4] ), .out(n1801) );
  xor2 U1357 ( .a(n1803), .b(n1799), .out(n1802) );
  xor2 U1358 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[1][2] ), .b(
        \mat_kron/mult_40_G2_G1_G1/ab[0][3] ), .out(n1804) );
  xor2 U1359 ( .a(n1806), .b(n1801), .out(n1805) );
  xor2 U1360 ( .a(n1808), .b(n1092), .out(n1807) );
  xor2 U1361 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[1][1] ), .b(
        \mat_kron/mult_40_G2_G1_G1/ab[0][2] ), .out(n1809) );
  xor2 U1362 ( .a(n1811), .b(n1804), .out(n1810) );
  xor2 U1363 ( .a(n1813), .b(n1814), .out(n1812) );
  xor2 U1364 ( .a(n1815), .b(n1816), .out(\mat_kron/mult_40_G2_G1_G1/A1[5] )
         );
  xor2 U1365 ( .a(n1817), .b(n1812), .out(\mat_kron/mult_40_G2_G1_G1/A1[3] )
         );
  xor2 U1366 ( .a(n1818), .b(n1810), .out(\mat_kron/mult_40_G2_G1_G1/A1[1] )
         );
  xor2 U1367 ( .a(\mat_kron/mult_40_G2_G1/ab[1][5] ), .b(
        \mat_kron/mult_40_G2_G1/ab[0][6] ), .out(n1121) );
  xor2 U1368 ( .a(n1819), .b(n1121), .out(n1127) );
  xor2 U1369 ( .a(n1821), .b(\mat_kron/mult_40_G2_G1/ab[0][5] ), .out(n1820)
         );
  xor2 U1370 ( .a(\mat_kron/mult_40_G2_G1/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G1/ab[0][4] ), .out(n1822) );
  xor2 U1371 ( .a(n1824), .b(n1820), .out(n1823) );
  xor2 U1372 ( .a(\mat_kron/mult_40_G2_G1/ab[1][2] ), .b(
        \mat_kron/mult_40_G2_G1/ab[0][3] ), .out(n1825) );
  xor2 U1373 ( .a(n1827), .b(n1822), .out(n1826) );
  xor2 U1374 ( .a(n1829), .b(n1136), .out(n1828) );
  xor2 U1375 ( .a(\mat_kron/mult_40_G2_G1/ab[1][1] ), .b(
        \mat_kron/mult_40_G2_G1/ab[0][2] ), .out(n1830) );
  xor2 U1376 ( .a(n1832), .b(n1825), .out(n1831) );
  xor2 U1377 ( .a(n1834), .b(n1835), .out(n1833) );
  xor2 U1378 ( .a(n1836), .b(n1837), .out(\mat_kron/mult_40_G2_G1/A1[5] ) );
  xor2 U1379 ( .a(n1838), .b(n1833), .out(\mat_kron/mult_40_G2_G1/A1[3] ) );
  xor2 U1380 ( .a(n1839), .b(n1831), .out(\mat_kron/mult_40_G2_G1/A1[1] ) );
  xor2 U1381 ( .a(\mat_kron/mult_40_G2/ab[1][5] ), .b(
        \mat_kron/mult_40_G2/ab[0][6] ), .out(n1165) );
  xor2 U1382 ( .a(n1840), .b(n1165), .out(n1171) );
  xor2 U1383 ( .a(n1842), .b(\mat_kron/mult_40_G2/ab[0][5] ), .out(n1841) );
  xor2 U1384 ( .a(\mat_kron/mult_40_G2/ab[1][3] ), .b(
        \mat_kron/mult_40_G2/ab[0][4] ), .out(n1843) );
  xor2 U1385 ( .a(n1845), .b(n1841), .out(n1844) );
  xor2 U1386 ( .a(\mat_kron/mult_40_G2/ab[1][2] ), .b(
        \mat_kron/mult_40_G2/ab[0][3] ), .out(n1846) );
  xor2 U1387 ( .a(n1848), .b(n1843), .out(n1847) );
  xor2 U1388 ( .a(n1850), .b(n1180), .out(n1849) );
  xor2 U1389 ( .a(\mat_kron/mult_40_G2/ab[1][1] ), .b(
        \mat_kron/mult_40_G2/ab[0][2] ), .out(n1851) );
  xor2 U1390 ( .a(n1853), .b(n1846), .out(n1852) );
  xor2 U1391 ( .a(n1855), .b(n1856), .out(n1854) );
  xor2 U1392 ( .a(n1857), .b(n1858), .out(\mat_kron/mult_40_G2/A1[5] ) );
  xor2 U1393 ( .a(n1859), .b(n1854), .out(\mat_kron/mult_40_G2/A1[3] ) );
  xor2 U1394 ( .a(n1860), .b(n1852), .out(\mat_kron/mult_40_G2/A1[1] ) );
  xor2 U1395 ( .a(\mat_kron/mult_40/ab[1][5] ), .b(\mat_kron/mult_40/ab[0][6] ), .out(n1209) );
  xor2 U1396 ( .a(n1861), .b(n1209), .out(n1215) );
  xor2 U1397 ( .a(n1863), .b(\mat_kron/mult_40/ab[0][5] ), .out(n1862) );
  xor2 U1398 ( .a(\mat_kron/mult_40/ab[1][3] ), .b(\mat_kron/mult_40/ab[0][4] ), .out(n1864) );
  xor2 U1399 ( .a(n1866), .b(n1862), .out(n1865) );
  xor2 U1400 ( .a(\mat_kron/mult_40/ab[1][2] ), .b(\mat_kron/mult_40/ab[0][3] ), .out(n1867) );
  xor2 U1401 ( .a(n1869), .b(n1864), .out(n1868) );
  xor2 U1402 ( .a(n1871), .b(n1224), .out(n1870) );
  xor2 U1403 ( .a(\mat_kron/mult_40/ab[1][1] ), .b(\mat_kron/mult_40/ab[0][2] ), .out(n1872) );
  xor2 U1404 ( .a(n1874), .b(n1867), .out(n1873) );
  xor2 U1405 ( .a(n1876), .b(n1877), .out(n1875) );
  xor2 U1406 ( .a(n1878), .b(n1879), .out(\mat_kron/mult_40/A1[5] ) );
  xor2 U1407 ( .a(n1880), .b(n1875), .out(\mat_kron/mult_40/A1[3] ) );
  xor2 U1408 ( .a(n1881), .b(n1873), .out(\mat_kron/mult_40/A1[1] ) );
  xor2 U1409 ( .a(n1298), .b(n1882), .out(m_sub[9]) );
  xor2 U1410 ( .a(n1883), .b(n1264), .out(m_sub[7]) );
  xor2 U1411 ( .a(n1884), .b(n1266), .out(m_sub[6]) );
  xor2 U1412 ( .a(n1885), .b(n1263), .out(m_sub[5]) );
  xor2 U1413 ( .a(n1886), .b(n1260), .out(m_sub[4]) );
  xor2 U1414 ( .a(n1887), .b(n1258), .out(m_sub[3]) );
  xor2 U1415 ( .a(n1888), .b(n1279), .out(m_sub[31]) );
  xor2 U1416 ( .a(n1889), .b(n1281), .out(m_sub[30]) );
  xor2 U1417 ( .a(n1890), .b(n1255), .out(m_sub[2]) );
  xor2 U1418 ( .a(n1891), .b(n1278), .out(m_sub[29]) );
  xor2 U1419 ( .a(n1892), .b(n1275), .out(m_sub[28]) );
  xor2 U1420 ( .a(n1893), .b(n1273), .out(m_sub[27]) );
  xor2 U1421 ( .a(n1894), .b(n1270), .out(m_sub[26]) );
  xor2 U1422 ( .a(n1268), .b(n1895), .out(m_sub[25]) );
  xor2 U1423 ( .a(n1896), .b(n1294), .out(m_sub[23]) );
  xor2 U1424 ( .a(n1897), .b(n1296), .out(m_sub[22]) );
  xor2 U1425 ( .a(n1898), .b(n1293), .out(m_sub[21]) );
  xor2 U1426 ( .a(n1899), .b(n1290), .out(m_sub[20]) );
  xor2 U1427 ( .a(n1253), .b(n1900), .out(m_sub[1]) );
  xor2 U1428 ( .a(n1901), .b(n1288), .out(m_sub[19]) );
  xor2 U1429 ( .a(n1902), .b(n1285), .out(m_sub[18]) );
  xor2 U1430 ( .a(n1283), .b(n1903), .out(m_sub[17]) );
  xor2 U1431 ( .a(n1904), .b(n1311), .out(m_sub[15]) );
  xor2 U1432 ( .a(n1905), .b(n1313), .out(m_sub[14]) );
  xor2 U1433 ( .a(n1906), .b(n1310), .out(m_sub[13]) );
  xor2 U1434 ( .a(n1907), .b(n1307), .out(m_sub[12]) );
  xor2 U1435 ( .a(n1908), .b(n1304), .out(m_sub[11]) );
  xor2 U1436 ( .a(n1909), .b(n1301), .out(m_sub[10]) );
  xor2 U1437 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[1][0] ), .b(
        \mat_mul/mult_37_G2_G1_G2/ab[0][1] ), .out(n1340) );
  xor2 U1438 ( .a(\mat_mul/mult_37_G2/ab[1][0] ), .b(
        \mat_mul/mult_37_G2/ab[0][1] ), .out(n1339) );
  xor2 U1439 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[1][0] ), .b(
        \mat_mul/mult_37_G2_G2_G2/ab[0][1] ), .out(n1316) );
  xor2 U1440 ( .a(\mat_mul/mult_37_G2_G2/ab[1][0] ), .b(
        \mat_mul/mult_37_G2_G2/ab[0][1] ), .out(n1315) );
  xor2 U1441 ( .a(n1911), .b(n1912), .out(n1910) );
  xor2 U1442 ( .a(n1913), .b(n1914), .out(m_mul[6]) );
  xor2 U1443 ( .a(n1915), .b(n1916), .out(m_mul[5]) );
  xor2 U1444 ( .a(n1917), .b(n1918), .out(m_mul[4]) );
  xor2 U1445 ( .a(n1919), .b(n1920), .out(m_mul[3]) );
  xor2 U1446 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[1][0] ), .b(
        \mat_mul/mult_37_G2_G1_G1/ab[0][1] ), .out(n1324) );
  xor2 U1447 ( .a(\mat_mul/mult_37/ab[1][0] ), .b(\mat_mul/mult_37/ab[0][1] ), 
        .out(n1323) );
  xor2 U1448 ( .a(n1922), .b(n1923), .out(n1921) );
  xor2 U1449 ( .a(n1924), .b(n1925), .out(m_mul[30]) );
  xor2 U1450 ( .a(n1926), .b(n1927), .out(m_mul[2]) );
  xor2 U1451 ( .a(n1928), .b(n1929), .out(m_mul[29]) );
  xor2 U1452 ( .a(n1930), .b(n1931), .out(m_mul[28]) );
  xor2 U1453 ( .a(n1932), .b(n1933), .out(m_mul[27]) );
  xor2 U1454 ( .a(n1934), .b(n1935), .out(m_mul[26]) );
  xor2 U1455 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[1][0] ), .b(
        \mat_mul/mult_37_G2_G2_G1/ab[0][1] ), .out(n1332) );
  xor2 U1456 ( .a(\mat_mul/mult_37_G2_G1/ab[1][0] ), .b(
        \mat_mul/mult_37_G2_G1/ab[0][1] ), .out(n1331) );
  xor2 U1457 ( .a(n1937), .b(n1938), .out(n1936) );
  xor2 U1458 ( .a(n1939), .b(n1940), .out(m_mul[22]) );
  xor2 U1459 ( .a(n1941), .b(n1942), .out(m_mul[21]) );
  xor2 U1460 ( .a(n1943), .b(n1944), .out(m_mul[20]) );
  xor2 U1461 ( .a(n1945), .b(n1946), .out(m_mul[19]) );
  xor2 U1462 ( .a(n1947), .b(n1948), .out(m_mul[18]) );
  xor2 U1463 ( .a(n1950), .b(n1951), .out(n1949) );
  xor2 U1464 ( .a(n1952), .b(n1953), .out(m_mul[14]) );
  xor2 U1465 ( .a(n1954), .b(n1955), .out(m_mul[13]) );
  xor2 U1466 ( .a(n1956), .b(n1957), .out(m_mul[12]) );
  xor2 U1467 ( .a(n1958), .b(n1959), .out(m_mul[11]) );
  xor2 U1468 ( .a(n1960), .b(n1961), .out(m_mul[10]) );
  xor2 U1469 ( .a(n1962), .b(n1351), .out(m_add[7]) );
  xor2 U1470 ( .a(n1353), .b(n1963), .out(m_add[6]) );
  xor2 U1471 ( .a(n1964), .b(n1965), .out(m_add[5]) );
  xor2 U1472 ( .a(n1966), .b(n1967), .out(m_add[4]) );
  xor2 U1473 ( .a(n1968), .b(n1969), .out(m_add[3]) );
  xor2 U1474 ( .a(n1970), .b(n1359), .out(m_add[31]) );
  xor2 U1475 ( .a(n1361), .b(n1971), .out(m_add[30]) );
  xor2 U1476 ( .a(n1972), .b(n1973), .out(m_add[2]) );
  xor2 U1477 ( .a(n1974), .b(n1975), .out(m_add[29]) );
  xor2 U1478 ( .a(n1976), .b(n1977), .out(m_add[28]) );
  xor2 U1479 ( .a(n1978), .b(n1979), .out(m_add[27]) );
  xor2 U1480 ( .a(n1980), .b(n1981), .out(m_add[26]) );
  xor2 U1481 ( .a(n1982), .b(n1367), .out(m_add[23]) );
  xor2 U1482 ( .a(n1369), .b(n1983), .out(m_add[22]) );
  xor2 U1483 ( .a(n1984), .b(n1985), .out(m_add[21]) );
  xor2 U1484 ( .a(n1986), .b(n1987), .out(m_add[20]) );
  xor2 U1485 ( .a(n1988), .b(n1989), .out(m_add[19]) );
  xor2 U1486 ( .a(n1990), .b(n1991), .out(m_add[18]) );
  xor2 U1487 ( .a(n1992), .b(n1375), .out(m_add[15]) );
  xor2 U1488 ( .a(n1377), .b(n1993), .out(m_add[14]) );
  xor2 U1489 ( .a(n1994), .b(n1995), .out(m_add[13]) );
  xor2 U1490 ( .a(n1996), .b(n1997), .out(m_add[12]) );
  xor2 U1491 ( .a(n1998), .b(n1999), .out(m_add[11]) );
  xor2 U1492 ( .a(n2000), .b(n2001), .out(m_add[10]) );
  nand2 U1493 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[0][3] ), .b(
        \mat_mul/mult_37_G2_G2_G2/ab[1][2] ), .out(n2002) );
  aoi22 U1494 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[2][2] ), .b(n207), .c(n2003), 
        .d(n1381), .out(n210) );
  nand2 U1495 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[1][3] ), .b(
        \mat_mul/mult_37_G2_G2_G2/ab[0][4] ), .out(n2004) );
  inv U1496 ( .in(\mat_mul/mult_37_G2_G2_G2/ab[2][3] ), .out(n2005) );
  aoi22 U1497 ( .a(n2007), .b(\mat_mul/mult_37_G2_G2_G2/ab[3][2] ), .c(n208), 
        .d(n1382), .out(n2006) );
  nand2 U1498 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[1][4] ), .b(
        \mat_mul/mult_37_G2_G2_G2/ab[0][5] ), .out(n2008) );
  oai22 U1499 ( .a(n2004), .b(n2005), .c(n200), .d(n1379), .out(n205) );
  nand2 U1500 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[0][2] ), .b(
        \mat_mul/mult_37_G2_G2_G2/ab[1][1] ), .out(n217) );
  aoi22 U1501 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[2][1] ), .b(n2010), .c(n215), 
        .d(n1384), .out(n2009) );
  oai22 U1502 ( .a(n2009), .b(n2011), .c(n218), .d(n1385), .out(n221) );
  inv U1503 ( .in(\mat_mul/mult_37_G2_G2_G2/ab[4][1] ), .out(n2012) );
  oai22 U1504 ( .a(n2013), .b(n2012), .c(n220), .d(n1394), .out(n223) );
  inv U1505 ( .in(\mat_mul/mult_37_G2_G2_G2/ab[5][1] ), .out(n2014) );
  nand2 U1506 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[0][1] ), .b(
        \mat_mul/mult_37_G2_G2_G2/ab[1][0] ), .out(n226) );
  aoi22 U1507 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[2][0] ), .b(n2015), .c(n224), 
        .d(n1389), .out(n229) );
  aoi22 U1508 ( .a(n2016), .b(\mat_mul/mult_37_G2_G2_G2/ab[3][0] ), .c(n227), 
        .d(n1390), .out(n232) );
  inv U1509 ( .in(\mat_mul/mult_37_G2_G2_G2/ab[4][0] ), .out(n231) );
  oai22 U1510 ( .a(n232), .b(n231), .c(n2017), .d(n2018), .out(n234) );
  aoi22 U1511 ( .a(n234), .b(\mat_mul/mult_37_G2_G2_G2/ab[5][0] ), .c(n2019), 
        .d(n1392), .out(n239) );
  nand2 U1512 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[0][3] ), .b(
        \mat_mul/mult_37_G2_G2_G1/ab[1][2] ), .out(n2020) );
  aoi22 U1513 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[2][2] ), .b(n251), .c(n2021), 
        .d(n1402), .out(n254) );
  nand2 U1514 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[1][3] ), .b(
        \mat_mul/mult_37_G2_G2_G1/ab[0][4] ), .out(n2022) );
  inv U1515 ( .in(\mat_mul/mult_37_G2_G2_G1/ab[2][3] ), .out(n2023) );
  aoi22 U1516 ( .a(n2025), .b(\mat_mul/mult_37_G2_G2_G1/ab[3][2] ), .c(n252), 
        .d(n1403), .out(n2024) );
  nand2 U1517 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[1][4] ), .b(
        \mat_mul/mult_37_G2_G2_G1/ab[0][5] ), .out(n2026) );
  oai22 U1518 ( .a(n2022), .b(n2023), .c(n244), .d(n1400), .out(n249) );
  nand2 U1519 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[0][2] ), .b(
        \mat_mul/mult_37_G2_G2_G1/ab[1][1] ), .out(n261) );
  aoi22 U1520 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[2][1] ), .b(n2028), .c(n259), 
        .d(n1405), .out(n2027) );
  oai22 U1521 ( .a(n2027), .b(n2029), .c(n262), .d(n1406), .out(n265) );
  inv U1522 ( .in(\mat_mul/mult_37_G2_G2_G1/ab[4][1] ), .out(n2030) );
  oai22 U1523 ( .a(n2031), .b(n2030), .c(n264), .d(n1415), .out(n267) );
  inv U1524 ( .in(\mat_mul/mult_37_G2_G2_G1/ab[5][1] ), .out(n2032) );
  nand2 U1525 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[0][1] ), .b(
        \mat_mul/mult_37_G2_G2_G1/ab[1][0] ), .out(n270) );
  aoi22 U1526 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[2][0] ), .b(n2033), .c(n268), 
        .d(n1410), .out(n273) );
  aoi22 U1527 ( .a(n2034), .b(\mat_mul/mult_37_G2_G2_G1/ab[3][0] ), .c(n271), 
        .d(n1411), .out(n276) );
  inv U1528 ( .in(\mat_mul/mult_37_G2_G2_G1/ab[4][0] ), .out(n275) );
  oai22 U1529 ( .a(n276), .b(n275), .c(n2035), .d(n2036), .out(n278) );
  aoi22 U1530 ( .a(n278), .b(\mat_mul/mult_37_G2_G2_G1/ab[5][0] ), .c(n2037), 
        .d(n1413), .out(n283) );
  nand2 U1531 ( .a(\mat_mul/mult_37_G2_G2/ab[0][3] ), .b(
        \mat_mul/mult_37_G2_G2/ab[1][2] ), .out(n2038) );
  aoi22 U1532 ( .a(\mat_mul/mult_37_G2_G2/ab[2][2] ), .b(n295), .c(n2039), .d(
        n1423), .out(n298) );
  nand2 U1533 ( .a(\mat_mul/mult_37_G2_G2/ab[1][3] ), .b(
        \mat_mul/mult_37_G2_G2/ab[0][4] ), .out(n2040) );
  inv U1534 ( .in(\mat_mul/mult_37_G2_G2/ab[2][3] ), .out(n2041) );
  aoi22 U1535 ( .a(n2043), .b(\mat_mul/mult_37_G2_G2/ab[3][2] ), .c(n296), .d(
        n1424), .out(n2042) );
  nand2 U1536 ( .a(\mat_mul/mult_37_G2_G2/ab[1][4] ), .b(
        \mat_mul/mult_37_G2_G2/ab[0][5] ), .out(n2044) );
  oai22 U1537 ( .a(n2040), .b(n2041), .c(n288), .d(n1421), .out(n293) );
  nand2 U1538 ( .a(\mat_mul/mult_37_G2_G2/ab[0][2] ), .b(
        \mat_mul/mult_37_G2_G2/ab[1][1] ), .out(n305) );
  aoi22 U1539 ( .a(\mat_mul/mult_37_G2_G2/ab[2][1] ), .b(n2046), .c(n303), .d(
        n1426), .out(n2045) );
  oai22 U1540 ( .a(n2045), .b(n2047), .c(n306), .d(n1427), .out(n309) );
  inv U1541 ( .in(\mat_mul/mult_37_G2_G2/ab[4][1] ), .out(n2048) );
  oai22 U1542 ( .a(n2049), .b(n2048), .c(n308), .d(n1436), .out(n311) );
  inv U1543 ( .in(\mat_mul/mult_37_G2_G2/ab[5][1] ), .out(n2050) );
  nand2 U1544 ( .a(\mat_mul/mult_37_G2_G2/ab[0][1] ), .b(
        \mat_mul/mult_37_G2_G2/ab[1][0] ), .out(n314) );
  aoi22 U1545 ( .a(\mat_mul/mult_37_G2_G2/ab[2][0] ), .b(n2051), .c(n312), .d(
        n1431), .out(n317) );
  aoi22 U1546 ( .a(n2052), .b(\mat_mul/mult_37_G2_G2/ab[3][0] ), .c(n315), .d(
        n1432), .out(n320) );
  inv U1547 ( .in(\mat_mul/mult_37_G2_G2/ab[4][0] ), .out(n319) );
  oai22 U1548 ( .a(n320), .b(n319), .c(n2053), .d(n2054), .out(n322) );
  aoi22 U1549 ( .a(n322), .b(\mat_mul/mult_37_G2_G2/ab[5][0] ), .c(n2055), .d(
        n1434), .out(n327) );
  nand2 U1550 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[0][3] ), .b(
        \mat_mul/mult_37_G2_G1_G2/ab[1][2] ), .out(n2056) );
  aoi22 U1551 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[2][2] ), .b(n339), .c(n2057), 
        .d(n1444), .out(n342) );
  nand2 U1552 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[1][3] ), .b(
        \mat_mul/mult_37_G2_G1_G2/ab[0][4] ), .out(n2058) );
  inv U1553 ( .in(\mat_mul/mult_37_G2_G1_G2/ab[2][3] ), .out(n2059) );
  aoi22 U1554 ( .a(n2061), .b(\mat_mul/mult_37_G2_G1_G2/ab[3][2] ), .c(n340), 
        .d(n1445), .out(n2060) );
  nand2 U1555 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[1][4] ), .b(
        \mat_mul/mult_37_G2_G1_G2/ab[0][5] ), .out(n2062) );
  oai22 U1556 ( .a(n2058), .b(n2059), .c(n332), .d(n1442), .out(n337) );
  nand2 U1557 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[0][2] ), .b(
        \mat_mul/mult_37_G2_G1_G2/ab[1][1] ), .out(n349) );
  aoi22 U1558 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[2][1] ), .b(n2064), .c(n347), 
        .d(n1447), .out(n2063) );
  oai22 U1559 ( .a(n2063), .b(n2065), .c(n350), .d(n1448), .out(n353) );
  inv U1560 ( .in(\mat_mul/mult_37_G2_G1_G2/ab[4][1] ), .out(n2066) );
  oai22 U1561 ( .a(n2067), .b(n2066), .c(n352), .d(n1457), .out(n355) );
  inv U1562 ( .in(\mat_mul/mult_37_G2_G1_G2/ab[5][1] ), .out(n2068) );
  nand2 U1563 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[0][1] ), .b(
        \mat_mul/mult_37_G2_G1_G2/ab[1][0] ), .out(n358) );
  aoi22 U1564 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[2][0] ), .b(n2069), .c(n356), 
        .d(n1452), .out(n361) );
  aoi22 U1565 ( .a(n2070), .b(\mat_mul/mult_37_G2_G1_G2/ab[3][0] ), .c(n359), 
        .d(n1453), .out(n364) );
  inv U1566 ( .in(\mat_mul/mult_37_G2_G1_G2/ab[4][0] ), .out(n363) );
  oai22 U1567 ( .a(n364), .b(n363), .c(n2071), .d(n2072), .out(n366) );
  aoi22 U1568 ( .a(n366), .b(\mat_mul/mult_37_G2_G1_G2/ab[5][0] ), .c(n2073), 
        .d(n1455), .out(n371) );
  nand2 U1569 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[0][3] ), .b(
        \mat_mul/mult_37_G2_G1_G1/ab[1][2] ), .out(n2074) );
  aoi22 U1570 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[2][2] ), .b(n383), .c(n2075), 
        .d(n1465), .out(n386) );
  nand2 U1571 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[1][3] ), .b(
        \mat_mul/mult_37_G2_G1_G1/ab[0][4] ), .out(n2076) );
  inv U1572 ( .in(\mat_mul/mult_37_G2_G1_G1/ab[2][3] ), .out(n2077) );
  aoi22 U1573 ( .a(n2079), .b(\mat_mul/mult_37_G2_G1_G1/ab[3][2] ), .c(n384), 
        .d(n1466), .out(n2078) );
  nand2 U1574 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[1][4] ), .b(
        \mat_mul/mult_37_G2_G1_G1/ab[0][5] ), .out(n2080) );
  oai22 U1575 ( .a(n2076), .b(n2077), .c(n376), .d(n1463), .out(n381) );
  nand2 U1576 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[0][2] ), .b(
        \mat_mul/mult_37_G2_G1_G1/ab[1][1] ), .out(n393) );
  aoi22 U1577 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[2][1] ), .b(n2082), .c(n391), 
        .d(n1468), .out(n2081) );
  oai22 U1578 ( .a(n2081), .b(n2083), .c(n394), .d(n1469), .out(n397) );
  inv U1579 ( .in(\mat_mul/mult_37_G2_G1_G1/ab[4][1] ), .out(n2084) );
  oai22 U1580 ( .a(n2085), .b(n2084), .c(n396), .d(n1478), .out(n399) );
  inv U1581 ( .in(\mat_mul/mult_37_G2_G1_G1/ab[5][1] ), .out(n2086) );
  nand2 U1582 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[0][1] ), .b(
        \mat_mul/mult_37_G2_G1_G1/ab[1][0] ), .out(n402) );
  aoi22 U1583 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[2][0] ), .b(n2087), .c(n400), 
        .d(n1473), .out(n405) );
  aoi22 U1584 ( .a(n2088), .b(\mat_mul/mult_37_G2_G1_G1/ab[3][0] ), .c(n403), 
        .d(n1474), .out(n408) );
  inv U1585 ( .in(\mat_mul/mult_37_G2_G1_G1/ab[4][0] ), .out(n407) );
  oai22 U1586 ( .a(n408), .b(n407), .c(n2089), .d(n2090), .out(n410) );
  aoi22 U1587 ( .a(n410), .b(\mat_mul/mult_37_G2_G1_G1/ab[5][0] ), .c(n2091), 
        .d(n1476), .out(n415) );
  nand2 U1588 ( .a(\mat_mul/mult_37_G2_G1/ab[0][3] ), .b(
        \mat_mul/mult_37_G2_G1/ab[1][2] ), .out(n2092) );
  aoi22 U1589 ( .a(\mat_mul/mult_37_G2_G1/ab[2][2] ), .b(n427), .c(n2093), .d(
        n1486), .out(n430) );
  nand2 U1590 ( .a(\mat_mul/mult_37_G2_G1/ab[1][3] ), .b(
        \mat_mul/mult_37_G2_G1/ab[0][4] ), .out(n2094) );
  inv U1591 ( .in(\mat_mul/mult_37_G2_G1/ab[2][3] ), .out(n2095) );
  aoi22 U1592 ( .a(n2097), .b(\mat_mul/mult_37_G2_G1/ab[3][2] ), .c(n428), .d(
        n1487), .out(n2096) );
  nand2 U1593 ( .a(\mat_mul/mult_37_G2_G1/ab[1][4] ), .b(
        \mat_mul/mult_37_G2_G1/ab[0][5] ), .out(n2098) );
  oai22 U1594 ( .a(n2094), .b(n2095), .c(n420), .d(n1484), .out(n425) );
  nand2 U1595 ( .a(\mat_mul/mult_37_G2_G1/ab[0][2] ), .b(
        \mat_mul/mult_37_G2_G1/ab[1][1] ), .out(n437) );
  aoi22 U1596 ( .a(\mat_mul/mult_37_G2_G1/ab[2][1] ), .b(n2100), .c(n435), .d(
        n1489), .out(n2099) );
  oai22 U1597 ( .a(n2099), .b(n2101), .c(n438), .d(n1490), .out(n441) );
  inv U1598 ( .in(\mat_mul/mult_37_G2_G1/ab[4][1] ), .out(n2102) );
  oai22 U1599 ( .a(n2103), .b(n2102), .c(n440), .d(n1499), .out(n443) );
  inv U1600 ( .in(\mat_mul/mult_37_G2_G1/ab[5][1] ), .out(n2104) );
  nand2 U1601 ( .a(\mat_mul/mult_37_G2_G1/ab[0][1] ), .b(
        \mat_mul/mult_37_G2_G1/ab[1][0] ), .out(n446) );
  aoi22 U1602 ( .a(\mat_mul/mult_37_G2_G1/ab[2][0] ), .b(n2105), .c(n444), .d(
        n1494), .out(n449) );
  aoi22 U1603 ( .a(n2106), .b(\mat_mul/mult_37_G2_G1/ab[3][0] ), .c(n447), .d(
        n1495), .out(n452) );
  inv U1604 ( .in(\mat_mul/mult_37_G2_G1/ab[4][0] ), .out(n451) );
  oai22 U1605 ( .a(n452), .b(n451), .c(n2107), .d(n2108), .out(n454) );
  aoi22 U1606 ( .a(n454), .b(\mat_mul/mult_37_G2_G1/ab[5][0] ), .c(n2109), .d(
        n1497), .out(n459) );
  nand2 U1607 ( .a(\mat_mul/mult_37_G2/ab[0][3] ), .b(
        \mat_mul/mult_37_G2/ab[1][2] ), .out(n2110) );
  aoi22 U1608 ( .a(\mat_mul/mult_37_G2/ab[2][2] ), .b(n471), .c(n2111), .d(
        n1507), .out(n474) );
  nand2 U1609 ( .a(\mat_mul/mult_37_G2/ab[1][3] ), .b(
        \mat_mul/mult_37_G2/ab[0][4] ), .out(n2112) );
  inv U1610 ( .in(\mat_mul/mult_37_G2/ab[2][3] ), .out(n2113) );
  aoi22 U1611 ( .a(n2115), .b(\mat_mul/mult_37_G2/ab[3][2] ), .c(n472), .d(
        n1508), .out(n2114) );
  nand2 U1612 ( .a(\mat_mul/mult_37_G2/ab[1][4] ), .b(
        \mat_mul/mult_37_G2/ab[0][5] ), .out(n2116) );
  oai22 U1613 ( .a(n2112), .b(n2113), .c(n464), .d(n1505), .out(n469) );
  nand2 U1614 ( .a(\mat_mul/mult_37_G2/ab[0][2] ), .b(
        \mat_mul/mult_37_G2/ab[1][1] ), .out(n481) );
  aoi22 U1615 ( .a(\mat_mul/mult_37_G2/ab[2][1] ), .b(n2118), .c(n479), .d(
        n1510), .out(n2117) );
  oai22 U1616 ( .a(n2117), .b(n2119), .c(n482), .d(n1511), .out(n485) );
  inv U1617 ( .in(\mat_mul/mult_37_G2/ab[4][1] ), .out(n2120) );
  oai22 U1618 ( .a(n2121), .b(n2120), .c(n484), .d(n1520), .out(n487) );
  inv U1619 ( .in(\mat_mul/mult_37_G2/ab[5][1] ), .out(n2122) );
  nand2 U1620 ( .a(\mat_mul/mult_37_G2/ab[0][1] ), .b(
        \mat_mul/mult_37_G2/ab[1][0] ), .out(n490) );
  aoi22 U1621 ( .a(\mat_mul/mult_37_G2/ab[2][0] ), .b(n2123), .c(n488), .d(
        n1515), .out(n493) );
  aoi22 U1622 ( .a(n2124), .b(\mat_mul/mult_37_G2/ab[3][0] ), .c(n491), .d(
        n1516), .out(n496) );
  inv U1623 ( .in(\mat_mul/mult_37_G2/ab[4][0] ), .out(n495) );
  oai22 U1624 ( .a(n496), .b(n495), .c(n2125), .d(n2126), .out(n498) );
  aoi22 U1625 ( .a(n498), .b(\mat_mul/mult_37_G2/ab[5][0] ), .c(n2127), .d(
        n1518), .out(n503) );
  nand2 U1626 ( .a(\mat_mul/mult_37/ab[0][3] ), .b(\mat_mul/mult_37/ab[1][2] ), 
        .out(n2128) );
  aoi22 U1627 ( .a(\mat_mul/mult_37/ab[2][2] ), .b(n515), .c(n2129), .d(n1528), 
        .out(n518) );
  nand2 U1628 ( .a(\mat_mul/mult_37/ab[1][3] ), .b(\mat_mul/mult_37/ab[0][4] ), 
        .out(n2130) );
  inv U1629 ( .in(\mat_mul/mult_37/ab[2][3] ), .out(n2131) );
  aoi22 U1630 ( .a(n2133), .b(\mat_mul/mult_37/ab[3][2] ), .c(n516), .d(n1529), 
        .out(n2132) );
  nand2 U1631 ( .a(\mat_mul/mult_37/ab[1][4] ), .b(\mat_mul/mult_37/ab[0][5] ), 
        .out(n2134) );
  oai22 U1632 ( .a(n2130), .b(n2131), .c(n508), .d(n1526), .out(n513) );
  nand2 U1633 ( .a(\mat_mul/mult_37/ab[0][2] ), .b(\mat_mul/mult_37/ab[1][1] ), 
        .out(n525) );
  aoi22 U1634 ( .a(\mat_mul/mult_37/ab[2][1] ), .b(n2136), .c(n523), .d(n1531), 
        .out(n2135) );
  oai22 U1635 ( .a(n2135), .b(n2137), .c(n526), .d(n1532), .out(n529) );
  inv U1636 ( .in(\mat_mul/mult_37/ab[4][1] ), .out(n2138) );
  oai22 U1637 ( .a(n2139), .b(n2138), .c(n528), .d(n1541), .out(n531) );
  inv U1638 ( .in(\mat_mul/mult_37/ab[5][1] ), .out(n2140) );
  nand2 U1639 ( .a(\mat_mul/mult_37/ab[0][1] ), .b(\mat_mul/mult_37/ab[1][0] ), 
        .out(n534) );
  aoi22 U1640 ( .a(\mat_mul/mult_37/ab[2][0] ), .b(n2141), .c(n532), .d(n1536), 
        .out(n537) );
  aoi22 U1641 ( .a(n2142), .b(\mat_mul/mult_37/ab[3][0] ), .c(n535), .d(n1537), 
        .out(n540) );
  inv U1642 ( .in(\mat_mul/mult_37/ab[4][0] ), .out(n539) );
  oai22 U1643 ( .a(n540), .b(n539), .c(n2143), .d(n2144), .out(n542) );
  aoi22 U1644 ( .a(n542), .b(\mat_mul/mult_37/ab[5][0] ), .c(n2145), .d(n1539), 
        .out(n547) );
  nand2 U1645 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[0][3] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[1][2] ), .out(n2146) );
  aoi22 U1646 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[2][2] ), .b(n559), .c(
        n2147), .d(n1549), .out(n562) );
  nand2 U1647 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[0][4] ), .out(n2148) );
  inv U1648 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/ab[2][3] ), .out(n2149) );
  aoi22 U1649 ( .a(n2151), .b(\mat_kron/mult_40_G2_G2_G2_G2/ab[3][2] ), .c(
        n560), .d(n1550), .out(n2150) );
  nand2 U1650 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[1][4] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[0][5] ), .out(n2152) );
  oai22 U1651 ( .a(n2148), .b(n2149), .c(n552), .d(n1547), .out(n557) );
  nand2 U1652 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[0][2] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[1][1] ), .out(n569) );
  aoi22 U1653 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[2][1] ), .b(n2154), .c(
        n567), .d(n1552), .out(n2153) );
  oai22 U1654 ( .a(n2153), .b(n2155), .c(n570), .d(n1553), .out(n573) );
  inv U1655 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/ab[4][1] ), .out(n2156) );
  oai22 U1656 ( .a(n2157), .b(n2156), .c(n572), .d(n1562), .out(n575) );
  inv U1657 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/ab[5][1] ), .out(n2158) );
  nand2 U1658 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[1][0] ), .out(n578) );
  aoi22 U1659 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[2][0] ), .b(n2159), .c(
        n576), .d(n1557), .out(n581) );
  aoi22 U1660 ( .a(n2160), .b(\mat_kron/mult_40_G2_G2_G2_G2/ab[3][0] ), .c(
        n579), .d(n1558), .out(n584) );
  inv U1661 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/ab[4][0] ), .out(n583) );
  oai22 U1662 ( .a(n584), .b(n583), .c(n2161), .d(n2162), .out(n586) );
  aoi22 U1663 ( .a(n586), .b(\mat_kron/mult_40_G2_G2_G2_G2/ab[5][0] ), .c(
        n2163), .d(n1560), .out(n591) );
  nand2 U1664 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[0][3] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[1][2] ), .out(n2164) );
  aoi22 U1665 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[2][2] ), .b(n603), .c(
        n2165), .d(n1570), .out(n606) );
  nand2 U1666 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[0][4] ), .out(n2166) );
  inv U1667 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/ab[2][3] ), .out(n2167) );
  aoi22 U1668 ( .a(n2169), .b(\mat_kron/mult_40_G2_G2_G2_G1/ab[3][2] ), .c(
        n604), .d(n1571), .out(n2168) );
  nand2 U1669 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[1][4] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[0][5] ), .out(n2170) );
  oai22 U1670 ( .a(n2166), .b(n2167), .c(n596), .d(n1568), .out(n601) );
  nand2 U1671 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[0][2] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[1][1] ), .out(n613) );
  aoi22 U1672 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[2][1] ), .b(n2172), .c(
        n611), .d(n1573), .out(n2171) );
  oai22 U1673 ( .a(n2171), .b(n2173), .c(n614), .d(n1574), .out(n617) );
  inv U1674 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/ab[4][1] ), .out(n2174) );
  oai22 U1675 ( .a(n2175), .b(n2174), .c(n616), .d(n1583), .out(n619) );
  inv U1676 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/ab[5][1] ), .out(n2176) );
  nand2 U1677 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[1][0] ), .out(n622) );
  aoi22 U1678 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[2][0] ), .b(n2177), .c(
        n620), .d(n1578), .out(n625) );
  aoi22 U1679 ( .a(n2178), .b(\mat_kron/mult_40_G2_G2_G2_G1/ab[3][0] ), .c(
        n623), .d(n1579), .out(n628) );
  inv U1680 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/ab[4][0] ), .out(n627) );
  oai22 U1681 ( .a(n628), .b(n627), .c(n2179), .d(n2180), .out(n630) );
  aoi22 U1682 ( .a(n630), .b(\mat_kron/mult_40_G2_G2_G2_G1/ab[5][0] ), .c(
        n2181), .d(n1581), .out(n635) );
  nand2 U1683 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[0][3] ), .b(
        \mat_kron/mult_40_G2_G2_G2/ab[1][2] ), .out(n2182) );
  aoi22 U1684 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[2][2] ), .b(n647), .c(n2183), 
        .d(n1591), .out(n650) );
  nand2 U1685 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G2_G2/ab[0][4] ), .out(n2184) );
  inv U1686 ( .in(\mat_kron/mult_40_G2_G2_G2/ab[2][3] ), .out(n2185) );
  aoi22 U1687 ( .a(n2187), .b(\mat_kron/mult_40_G2_G2_G2/ab[3][2] ), .c(n648), 
        .d(n1592), .out(n2186) );
  nand2 U1688 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[1][4] ), .b(
        \mat_kron/mult_40_G2_G2_G2/ab[0][5] ), .out(n2188) );
  oai22 U1689 ( .a(n2184), .b(n2185), .c(n640), .d(n1589), .out(n645) );
  nand2 U1690 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[0][2] ), .b(
        \mat_kron/mult_40_G2_G2_G2/ab[1][1] ), .out(n657) );
  aoi22 U1691 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[2][1] ), .b(n2190), .c(n655), 
        .d(n1594), .out(n2189) );
  oai22 U1692 ( .a(n2189), .b(n2191), .c(n658), .d(n1595), .out(n661) );
  inv U1693 ( .in(\mat_kron/mult_40_G2_G2_G2/ab[4][1] ), .out(n2192) );
  oai22 U1694 ( .a(n2193), .b(n2192), .c(n660), .d(n1604), .out(n663) );
  inv U1695 ( .in(\mat_kron/mult_40_G2_G2_G2/ab[5][1] ), .out(n2194) );
  nand2 U1696 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G2_G2/ab[1][0] ), .out(n666) );
  aoi22 U1697 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[2][0] ), .b(n2195), .c(n664), 
        .d(n1599), .out(n669) );
  aoi22 U1698 ( .a(n2196), .b(\mat_kron/mult_40_G2_G2_G2/ab[3][0] ), .c(n667), 
        .d(n1600), .out(n672) );
  inv U1699 ( .in(\mat_kron/mult_40_G2_G2_G2/ab[4][0] ), .out(n671) );
  oai22 U1700 ( .a(n672), .b(n671), .c(n2197), .d(n2198), .out(n674) );
  aoi22 U1701 ( .a(n674), .b(\mat_kron/mult_40_G2_G2_G2/ab[5][0] ), .c(n2199), 
        .d(n1602), .out(n679) );
  nand2 U1702 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[0][3] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[1][2] ), .out(n2200) );
  aoi22 U1703 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[2][2] ), .b(n691), .c(
        n2201), .d(n1612), .out(n694) );
  nand2 U1704 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[0][4] ), .out(n2202) );
  inv U1705 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/ab[2][3] ), .out(n2203) );
  aoi22 U1706 ( .a(n2205), .b(\mat_kron/mult_40_G2_G2_G1_G2/ab[3][2] ), .c(
        n692), .d(n1613), .out(n2204) );
  nand2 U1707 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[1][4] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[0][5] ), .out(n2206) );
  oai22 U1708 ( .a(n2202), .b(n2203), .c(n684), .d(n1610), .out(n689) );
  nand2 U1709 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[0][2] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[1][1] ), .out(n701) );
  aoi22 U1710 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[2][1] ), .b(n2208), .c(
        n699), .d(n1615), .out(n2207) );
  oai22 U1711 ( .a(n2207), .b(n2209), .c(n702), .d(n1616), .out(n705) );
  inv U1712 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/ab[4][1] ), .out(n2210) );
  oai22 U1713 ( .a(n2211), .b(n2210), .c(n704), .d(n1625), .out(n707) );
  inv U1714 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/ab[5][1] ), .out(n2212) );
  nand2 U1715 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[1][0] ), .out(n710) );
  aoi22 U1716 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[2][0] ), .b(n2213), .c(
        n708), .d(n1620), .out(n713) );
  aoi22 U1717 ( .a(n2214), .b(\mat_kron/mult_40_G2_G2_G1_G2/ab[3][0] ), .c(
        n711), .d(n1621), .out(n716) );
  inv U1718 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/ab[4][0] ), .out(n715) );
  oai22 U1719 ( .a(n716), .b(n715), .c(n2215), .d(n2216), .out(n718) );
  aoi22 U1720 ( .a(n718), .b(\mat_kron/mult_40_G2_G2_G1_G2/ab[5][0] ), .c(
        n2217), .d(n1623), .out(n723) );
  nand2 U1721 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[0][3] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[1][2] ), .out(n2218) );
  aoi22 U1722 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[2][2] ), .b(n735), .c(
        n2219), .d(n1633), .out(n738) );
  nand2 U1723 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[0][4] ), .out(n2220) );
  inv U1724 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/ab[2][3] ), .out(n2221) );
  aoi22 U1725 ( .a(n2223), .b(\mat_kron/mult_40_G2_G2_G1_G1/ab[3][2] ), .c(
        n736), .d(n1634), .out(n2222) );
  nand2 U1726 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[1][4] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[0][5] ), .out(n2224) );
  oai22 U1727 ( .a(n2220), .b(n2221), .c(n728), .d(n1631), .out(n733) );
  nand2 U1728 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[0][2] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[1][1] ), .out(n745) );
  aoi22 U1729 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[2][1] ), .b(n2226), .c(
        n743), .d(n1636), .out(n2225) );
  oai22 U1730 ( .a(n2225), .b(n2227), .c(n746), .d(n1637), .out(n749) );
  inv U1731 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/ab[4][1] ), .out(n2228) );
  oai22 U1732 ( .a(n2229), .b(n2228), .c(n748), .d(n1646), .out(n751) );
  inv U1733 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/ab[5][1] ), .out(n2230) );
  nand2 U1734 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[1][0] ), .out(n754) );
  aoi22 U1735 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[2][0] ), .b(n2231), .c(
        n752), .d(n1641), .out(n757) );
  aoi22 U1736 ( .a(n2232), .b(\mat_kron/mult_40_G2_G2_G1_G1/ab[3][0] ), .c(
        n755), .d(n1642), .out(n760) );
  inv U1737 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/ab[4][0] ), .out(n759) );
  oai22 U1738 ( .a(n760), .b(n759), .c(n2233), .d(n2234), .out(n762) );
  aoi22 U1739 ( .a(n762), .b(\mat_kron/mult_40_G2_G2_G1_G1/ab[5][0] ), .c(
        n2235), .d(n1644), .out(n767) );
  nand2 U1740 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[0][3] ), .b(
        \mat_kron/mult_40_G2_G2_G1/ab[1][2] ), .out(n2236) );
  aoi22 U1741 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[2][2] ), .b(n779), .c(n2237), 
        .d(n1654), .out(n782) );
  nand2 U1742 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G2_G1/ab[0][4] ), .out(n2238) );
  inv U1743 ( .in(\mat_kron/mult_40_G2_G2_G1/ab[2][3] ), .out(n2239) );
  aoi22 U1744 ( .a(n2241), .b(\mat_kron/mult_40_G2_G2_G1/ab[3][2] ), .c(n780), 
        .d(n1655), .out(n2240) );
  nand2 U1745 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[1][4] ), .b(
        \mat_kron/mult_40_G2_G2_G1/ab[0][5] ), .out(n2242) );
  oai22 U1746 ( .a(n2238), .b(n2239), .c(n772), .d(n1652), .out(n777) );
  nand2 U1747 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[0][2] ), .b(
        \mat_kron/mult_40_G2_G2_G1/ab[1][1] ), .out(n789) );
  aoi22 U1748 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[2][1] ), .b(n2244), .c(n787), 
        .d(n1657), .out(n2243) );
  oai22 U1749 ( .a(n2243), .b(n2245), .c(n790), .d(n1658), .out(n793) );
  inv U1750 ( .in(\mat_kron/mult_40_G2_G2_G1/ab[4][1] ), .out(n2246) );
  oai22 U1751 ( .a(n2247), .b(n2246), .c(n792), .d(n1667), .out(n795) );
  inv U1752 ( .in(\mat_kron/mult_40_G2_G2_G1/ab[5][1] ), .out(n2248) );
  nand2 U1753 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G2_G1/ab[1][0] ), .out(n798) );
  aoi22 U1754 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[2][0] ), .b(n2249), .c(n796), 
        .d(n1662), .out(n801) );
  aoi22 U1755 ( .a(n2250), .b(\mat_kron/mult_40_G2_G2_G1/ab[3][0] ), .c(n799), 
        .d(n1663), .out(n804) );
  inv U1756 ( .in(\mat_kron/mult_40_G2_G2_G1/ab[4][0] ), .out(n803) );
  oai22 U1757 ( .a(n804), .b(n803), .c(n2251), .d(n2252), .out(n806) );
  aoi22 U1758 ( .a(n806), .b(\mat_kron/mult_40_G2_G2_G1/ab[5][0] ), .c(n2253), 
        .d(n1665), .out(n811) );
  nand2 U1759 ( .a(\mat_kron/mult_40_G2_G2/ab[0][3] ), .b(
        \mat_kron/mult_40_G2_G2/ab[1][2] ), .out(n2254) );
  aoi22 U1760 ( .a(\mat_kron/mult_40_G2_G2/ab[2][2] ), .b(n823), .c(n2255), 
        .d(n1675), .out(n826) );
  nand2 U1761 ( .a(\mat_kron/mult_40_G2_G2/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G2/ab[0][4] ), .out(n2256) );
  inv U1762 ( .in(\mat_kron/mult_40_G2_G2/ab[2][3] ), .out(n2257) );
  aoi22 U1763 ( .a(n2259), .b(\mat_kron/mult_40_G2_G2/ab[3][2] ), .c(n824), 
        .d(n1676), .out(n2258) );
  nand2 U1764 ( .a(\mat_kron/mult_40_G2_G2/ab[1][4] ), .b(
        \mat_kron/mult_40_G2_G2/ab[0][5] ), .out(n2260) );
  oai22 U1765 ( .a(n2256), .b(n2257), .c(n816), .d(n1673), .out(n821) );
  nand2 U1766 ( .a(\mat_kron/mult_40_G2_G2/ab[0][2] ), .b(
        \mat_kron/mult_40_G2_G2/ab[1][1] ), .out(n833) );
  aoi22 U1767 ( .a(\mat_kron/mult_40_G2_G2/ab[2][1] ), .b(n2262), .c(n831), 
        .d(n1678), .out(n2261) );
  oai22 U1768 ( .a(n2261), .b(n2263), .c(n834), .d(n1679), .out(n837) );
  inv U1769 ( .in(\mat_kron/mult_40_G2_G2/ab[4][1] ), .out(n2264) );
  oai22 U1770 ( .a(n2265), .b(n2264), .c(n836), .d(n1688), .out(n839) );
  inv U1771 ( .in(\mat_kron/mult_40_G2_G2/ab[5][1] ), .out(n2266) );
  nand2 U1772 ( .a(\mat_kron/mult_40_G2_G2/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G2/ab[1][0] ), .out(n842) );
  aoi22 U1773 ( .a(\mat_kron/mult_40_G2_G2/ab[2][0] ), .b(n2267), .c(n840), 
        .d(n1683), .out(n845) );
  aoi22 U1774 ( .a(n2268), .b(\mat_kron/mult_40_G2_G2/ab[3][0] ), .c(n843), 
        .d(n1684), .out(n848) );
  inv U1775 ( .in(\mat_kron/mult_40_G2_G2/ab[4][0] ), .out(n847) );
  oai22 U1776 ( .a(n848), .b(n847), .c(n2269), .d(n2270), .out(n850) );
  aoi22 U1777 ( .a(n850), .b(\mat_kron/mult_40_G2_G2/ab[5][0] ), .c(n2271), 
        .d(n1686), .out(n855) );
  nand2 U1778 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[0][3] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[1][2] ), .out(n2272) );
  aoi22 U1779 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[2][2] ), .b(n867), .c(
        n2273), .d(n1696), .out(n870) );
  nand2 U1780 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[0][4] ), .out(n2274) );
  inv U1781 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/ab[2][3] ), .out(n2275) );
  aoi22 U1782 ( .a(n2277), .b(\mat_kron/mult_40_G2_G1_G2_G2/ab[3][2] ), .c(
        n868), .d(n1697), .out(n2276) );
  nand2 U1783 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[1][4] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[0][5] ), .out(n2278) );
  oai22 U1784 ( .a(n2274), .b(n2275), .c(n860), .d(n1694), .out(n865) );
  nand2 U1785 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[0][2] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[1][1] ), .out(n877) );
  aoi22 U1786 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[2][1] ), .b(n2280), .c(
        n875), .d(n1699), .out(n2279) );
  oai22 U1787 ( .a(n2279), .b(n2281), .c(n878), .d(n1700), .out(n881) );
  inv U1788 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/ab[4][1] ), .out(n2282) );
  oai22 U1789 ( .a(n2283), .b(n2282), .c(n880), .d(n1709), .out(n883) );
  inv U1790 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/ab[5][1] ), .out(n2284) );
  nand2 U1791 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[1][0] ), .out(n886) );
  aoi22 U1792 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[2][0] ), .b(n2285), .c(
        n884), .d(n1704), .out(n889) );
  aoi22 U1793 ( .a(n2286), .b(\mat_kron/mult_40_G2_G1_G2_G2/ab[3][0] ), .c(
        n887), .d(n1705), .out(n892) );
  inv U1794 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/ab[4][0] ), .out(n891) );
  oai22 U1795 ( .a(n892), .b(n891), .c(n2287), .d(n2288), .out(n894) );
  aoi22 U1796 ( .a(n894), .b(\mat_kron/mult_40_G2_G1_G2_G2/ab[5][0] ), .c(
        n2289), .d(n1707), .out(n899) );
  nand2 U1797 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[0][3] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[1][2] ), .out(n2290) );
  aoi22 U1798 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[2][2] ), .b(n911), .c(
        n2291), .d(n1717), .out(n914) );
  nand2 U1799 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[0][4] ), .out(n2292) );
  inv U1800 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/ab[2][3] ), .out(n2293) );
  aoi22 U1801 ( .a(n2295), .b(\mat_kron/mult_40_G2_G1_G2_G1/ab[3][2] ), .c(
        n912), .d(n1718), .out(n2294) );
  nand2 U1802 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[1][4] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[0][5] ), .out(n2296) );
  oai22 U1803 ( .a(n2292), .b(n2293), .c(n904), .d(n1715), .out(n909) );
  nand2 U1804 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[0][2] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[1][1] ), .out(n921) );
  aoi22 U1805 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[2][1] ), .b(n2298), .c(
        n919), .d(n1720), .out(n2297) );
  oai22 U1806 ( .a(n2297), .b(n2299), .c(n922), .d(n1721), .out(n925) );
  inv U1807 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/ab[4][1] ), .out(n2300) );
  oai22 U1808 ( .a(n2301), .b(n2300), .c(n924), .d(n1730), .out(n927) );
  inv U1809 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/ab[5][1] ), .out(n2302) );
  nand2 U1810 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[1][0] ), .out(n930) );
  aoi22 U1811 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[2][0] ), .b(n2303), .c(
        n928), .d(n1725), .out(n933) );
  aoi22 U1812 ( .a(n2304), .b(\mat_kron/mult_40_G2_G1_G2_G1/ab[3][0] ), .c(
        n931), .d(n1726), .out(n936) );
  inv U1813 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/ab[4][0] ), .out(n935) );
  oai22 U1814 ( .a(n936), .b(n935), .c(n2305), .d(n2306), .out(n938) );
  aoi22 U1815 ( .a(n938), .b(\mat_kron/mult_40_G2_G1_G2_G1/ab[5][0] ), .c(
        n2307), .d(n1728), .out(n943) );
  nand2 U1816 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[0][3] ), .b(
        \mat_kron/mult_40_G2_G1_G2/ab[1][2] ), .out(n2308) );
  aoi22 U1817 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[2][2] ), .b(n955), .c(n2309), 
        .d(n1738), .out(n958) );
  nand2 U1818 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G1_G2/ab[0][4] ), .out(n2310) );
  inv U1819 ( .in(\mat_kron/mult_40_G2_G1_G2/ab[2][3] ), .out(n2311) );
  aoi22 U1820 ( .a(n2313), .b(\mat_kron/mult_40_G2_G1_G2/ab[3][2] ), .c(n956), 
        .d(n1739), .out(n2312) );
  nand2 U1821 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[1][4] ), .b(
        \mat_kron/mult_40_G2_G1_G2/ab[0][5] ), .out(n2314) );
  oai22 U1822 ( .a(n2310), .b(n2311), .c(n948), .d(n1736), .out(n953) );
  nand2 U1823 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[0][2] ), .b(
        \mat_kron/mult_40_G2_G1_G2/ab[1][1] ), .out(n965) );
  aoi22 U1824 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[2][1] ), .b(n2316), .c(n963), 
        .d(n1741), .out(n2315) );
  oai22 U1825 ( .a(n2315), .b(n2317), .c(n966), .d(n1742), .out(n969) );
  inv U1826 ( .in(\mat_kron/mult_40_G2_G1_G2/ab[4][1] ), .out(n2318) );
  oai22 U1827 ( .a(n2319), .b(n2318), .c(n968), .d(n1751), .out(n971) );
  inv U1828 ( .in(\mat_kron/mult_40_G2_G1_G2/ab[5][1] ), .out(n2320) );
  nand2 U1829 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G1_G2/ab[1][0] ), .out(n974) );
  aoi22 U1830 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[2][0] ), .b(n2321), .c(n972), 
        .d(n1746), .out(n977) );
  aoi22 U1831 ( .a(n2322), .b(\mat_kron/mult_40_G2_G1_G2/ab[3][0] ), .c(n975), 
        .d(n1747), .out(n980) );
  inv U1832 ( .in(\mat_kron/mult_40_G2_G1_G2/ab[4][0] ), .out(n979) );
  oai22 U1833 ( .a(n980), .b(n979), .c(n2323), .d(n2324), .out(n982) );
  aoi22 U1834 ( .a(n982), .b(\mat_kron/mult_40_G2_G1_G2/ab[5][0] ), .c(n2325), 
        .d(n1749), .out(n987) );
  nand2 U1835 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[0][3] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[1][2] ), .out(n2326) );
  aoi22 U1836 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[2][2] ), .b(n999), .c(
        n2327), .d(n1759), .out(n1002) );
  nand2 U1837 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[0][4] ), .out(n2328) );
  inv U1838 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/ab[2][3] ), .out(n2329) );
  aoi22 U1839 ( .a(n2331), .b(\mat_kron/mult_40_G2_G1_G1_G2/ab[3][2] ), .c(
        n1000), .d(n1760), .out(n2330) );
  nand2 U1840 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[1][4] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[0][5] ), .out(n2332) );
  oai22 U1841 ( .a(n2328), .b(n2329), .c(n992), .d(n1757), .out(n997) );
  nand2 U1842 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[0][2] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[1][1] ), .out(n1009) );
  aoi22 U1843 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[2][1] ), .b(n2334), .c(
        n1007), .d(n1762), .out(n2333) );
  oai22 U1844 ( .a(n2333), .b(n2335), .c(n1010), .d(n1763), .out(n1013) );
  inv U1845 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/ab[4][1] ), .out(n2336) );
  oai22 U1846 ( .a(n2337), .b(n2336), .c(n1012), .d(n1772), .out(n1015) );
  inv U1847 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/ab[5][1] ), .out(n2338) );
  nand2 U1848 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[1][0] ), .out(n1018) );
  aoi22 U1849 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[2][0] ), .b(n2339), .c(
        n1016), .d(n1767), .out(n1021) );
  aoi22 U1850 ( .a(n2340), .b(\mat_kron/mult_40_G2_G1_G1_G2/ab[3][0] ), .c(
        n1019), .d(n1768), .out(n1024) );
  inv U1851 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/ab[4][0] ), .out(n1023) );
  oai22 U1852 ( .a(n1024), .b(n1023), .c(n2341), .d(n2342), .out(n1026) );
  aoi22 U1853 ( .a(n1026), .b(\mat_kron/mult_40_G2_G1_G1_G2/ab[5][0] ), .c(
        n2343), .d(n1770), .out(n1031) );
  nand2 U1854 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[0][3] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[1][2] ), .out(n2344) );
  aoi22 U1855 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[2][2] ), .b(n1043), .c(
        n2345), .d(n1780), .out(n1046) );
  nand2 U1856 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[0][4] ), .out(n2346) );
  inv U1857 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/ab[2][3] ), .out(n2347) );
  aoi22 U1858 ( .a(n2349), .b(\mat_kron/mult_40_G2_G1_G1_G1/ab[3][2] ), .c(
        n1044), .d(n1781), .out(n2348) );
  nand2 U1859 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[1][4] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[0][5] ), .out(n2350) );
  oai22 U1860 ( .a(n2346), .b(n2347), .c(n1036), .d(n1778), .out(n1041) );
  nand2 U1861 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[0][2] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[1][1] ), .out(n1053) );
  aoi22 U1862 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[2][1] ), .b(n2352), .c(
        n1051), .d(n1783), .out(n2351) );
  oai22 U1863 ( .a(n2351), .b(n2353), .c(n1054), .d(n1784), .out(n1057) );
  inv U1864 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/ab[4][1] ), .out(n2354) );
  oai22 U1865 ( .a(n2355), .b(n2354), .c(n1056), .d(n1793), .out(n1059) );
  inv U1866 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/ab[5][1] ), .out(n2356) );
  nand2 U1867 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[1][0] ), .out(n1062) );
  aoi22 U1868 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[2][0] ), .b(n2357), .c(
        n1060), .d(n1788), .out(n1065) );
  aoi22 U1869 ( .a(n2358), .b(\mat_kron/mult_40_G2_G1_G1_G1/ab[3][0] ), .c(
        n1063), .d(n1789), .out(n1068) );
  inv U1870 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/ab[4][0] ), .out(n1067) );
  oai22 U1871 ( .a(n1068), .b(n1067), .c(n2359), .d(n2360), .out(n1070) );
  aoi22 U1872 ( .a(n1070), .b(\mat_kron/mult_40_G2_G1_G1_G1/ab[5][0] ), .c(
        n2361), .d(n1791), .out(n1075) );
  nand2 U1873 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[0][3] ), .b(
        \mat_kron/mult_40_G2_G1_G1/ab[1][2] ), .out(n2362) );
  aoi22 U1874 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[2][2] ), .b(n1087), .c(n2363), 
        .d(n1801), .out(n1090) );
  nand2 U1875 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G1_G1/ab[0][4] ), .out(n2364) );
  inv U1876 ( .in(\mat_kron/mult_40_G2_G1_G1/ab[2][3] ), .out(n2365) );
  aoi22 U1877 ( .a(n2367), .b(\mat_kron/mult_40_G2_G1_G1/ab[3][2] ), .c(n1088), 
        .d(n1802), .out(n2366) );
  nand2 U1878 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[1][4] ), .b(
        \mat_kron/mult_40_G2_G1_G1/ab[0][5] ), .out(n2368) );
  oai22 U1879 ( .a(n2364), .b(n2365), .c(n1080), .d(n1799), .out(n1085) );
  nand2 U1880 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[0][2] ), .b(
        \mat_kron/mult_40_G2_G1_G1/ab[1][1] ), .out(n1097) );
  aoi22 U1881 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[2][1] ), .b(n2370), .c(n1095), 
        .d(n1804), .out(n2369) );
  oai22 U1882 ( .a(n2369), .b(n2371), .c(n1098), .d(n1805), .out(n1101) );
  inv U1883 ( .in(\mat_kron/mult_40_G2_G1_G1/ab[4][1] ), .out(n2372) );
  oai22 U1884 ( .a(n2373), .b(n2372), .c(n1100), .d(n1814), .out(n1103) );
  inv U1885 ( .in(\mat_kron/mult_40_G2_G1_G1/ab[5][1] ), .out(n2374) );
  nand2 U1886 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G1_G1/ab[1][0] ), .out(n1106) );
  aoi22 U1887 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[2][0] ), .b(n2375), .c(n1104), 
        .d(n1809), .out(n1109) );
  aoi22 U1888 ( .a(n2376), .b(\mat_kron/mult_40_G2_G1_G1/ab[3][0] ), .c(n1107), 
        .d(n1810), .out(n1112) );
  inv U1889 ( .in(\mat_kron/mult_40_G2_G1_G1/ab[4][0] ), .out(n1111) );
  oai22 U1890 ( .a(n1112), .b(n1111), .c(n2377), .d(n2378), .out(n1114) );
  aoi22 U1891 ( .a(n1114), .b(\mat_kron/mult_40_G2_G1_G1/ab[5][0] ), .c(n2379), 
        .d(n1812), .out(n1119) );
  nand2 U1892 ( .a(\mat_kron/mult_40_G2_G1/ab[0][3] ), .b(
        \mat_kron/mult_40_G2_G1/ab[1][2] ), .out(n2380) );
  aoi22 U1893 ( .a(\mat_kron/mult_40_G2_G1/ab[2][2] ), .b(n1131), .c(n2381), 
        .d(n1822), .out(n1134) );
  nand2 U1894 ( .a(\mat_kron/mult_40_G2_G1/ab[1][3] ), .b(
        \mat_kron/mult_40_G2_G1/ab[0][4] ), .out(n2382) );
  inv U1895 ( .in(\mat_kron/mult_40_G2_G1/ab[2][3] ), .out(n2383) );
  aoi22 U1896 ( .a(n2385), .b(\mat_kron/mult_40_G2_G1/ab[3][2] ), .c(n1132), 
        .d(n1823), .out(n2384) );
  nand2 U1897 ( .a(\mat_kron/mult_40_G2_G1/ab[1][4] ), .b(
        \mat_kron/mult_40_G2_G1/ab[0][5] ), .out(n2386) );
  oai22 U1898 ( .a(n2382), .b(n2383), .c(n1124), .d(n1820), .out(n1129) );
  nand2 U1899 ( .a(\mat_kron/mult_40_G2_G1/ab[0][2] ), .b(
        \mat_kron/mult_40_G2_G1/ab[1][1] ), .out(n1141) );
  aoi22 U1900 ( .a(\mat_kron/mult_40_G2_G1/ab[2][1] ), .b(n2388), .c(n1139), 
        .d(n1825), .out(n2387) );
  oai22 U1901 ( .a(n2387), .b(n2389), .c(n1142), .d(n1826), .out(n1145) );
  inv U1902 ( .in(\mat_kron/mult_40_G2_G1/ab[4][1] ), .out(n2390) );
  oai22 U1903 ( .a(n2391), .b(n2390), .c(n1144), .d(n1835), .out(n1147) );
  inv U1904 ( .in(\mat_kron/mult_40_G2_G1/ab[5][1] ), .out(n2392) );
  nand2 U1905 ( .a(\mat_kron/mult_40_G2_G1/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G1/ab[1][0] ), .out(n1150) );
  aoi22 U1906 ( .a(\mat_kron/mult_40_G2_G1/ab[2][0] ), .b(n2393), .c(n1148), 
        .d(n1830), .out(n1153) );
  aoi22 U1907 ( .a(n2394), .b(\mat_kron/mult_40_G2_G1/ab[3][0] ), .c(n1151), 
        .d(n1831), .out(n1156) );
  inv U1908 ( .in(\mat_kron/mult_40_G2_G1/ab[4][0] ), .out(n1155) );
  oai22 U1909 ( .a(n1156), .b(n1155), .c(n2395), .d(n2396), .out(n1158) );
  aoi22 U1910 ( .a(n1158), .b(\mat_kron/mult_40_G2_G1/ab[5][0] ), .c(n2397), 
        .d(n1833), .out(n1163) );
  nand2 U1911 ( .a(\mat_kron/mult_40_G2/ab[0][3] ), .b(
        \mat_kron/mult_40_G2/ab[1][2] ), .out(n2398) );
  aoi22 U1912 ( .a(\mat_kron/mult_40_G2/ab[2][2] ), .b(n1175), .c(n2399), .d(
        n1843), .out(n1178) );
  nand2 U1913 ( .a(\mat_kron/mult_40_G2/ab[1][3] ), .b(
        \mat_kron/mult_40_G2/ab[0][4] ), .out(n2400) );
  inv U1914 ( .in(\mat_kron/mult_40_G2/ab[2][3] ), .out(n2401) );
  aoi22 U1915 ( .a(n2403), .b(\mat_kron/mult_40_G2/ab[3][2] ), .c(n1176), .d(
        n1844), .out(n2402) );
  nand2 U1916 ( .a(\mat_kron/mult_40_G2/ab[1][4] ), .b(
        \mat_kron/mult_40_G2/ab[0][5] ), .out(n2404) );
  oai22 U1917 ( .a(n2400), .b(n2401), .c(n1168), .d(n1841), .out(n1173) );
  nand2 U1918 ( .a(\mat_kron/mult_40_G2/ab[0][2] ), .b(
        \mat_kron/mult_40_G2/ab[1][1] ), .out(n1185) );
  aoi22 U1919 ( .a(\mat_kron/mult_40_G2/ab[2][1] ), .b(n2406), .c(n1183), .d(
        n1846), .out(n2405) );
  oai22 U1920 ( .a(n2405), .b(n2407), .c(n1186), .d(n1847), .out(n1189) );
  inv U1921 ( .in(\mat_kron/mult_40_G2/ab[4][1] ), .out(n2408) );
  oai22 U1922 ( .a(n2409), .b(n2408), .c(n1188), .d(n1856), .out(n1191) );
  inv U1923 ( .in(\mat_kron/mult_40_G2/ab[5][1] ), .out(n2410) );
  nand2 U1924 ( .a(\mat_kron/mult_40_G2/ab[0][1] ), .b(
        \mat_kron/mult_40_G2/ab[1][0] ), .out(n1194) );
  aoi22 U1925 ( .a(\mat_kron/mult_40_G2/ab[2][0] ), .b(n2411), .c(n1192), .d(
        n1851), .out(n1197) );
  aoi22 U1926 ( .a(n2412), .b(\mat_kron/mult_40_G2/ab[3][0] ), .c(n1195), .d(
        n1852), .out(n1200) );
  inv U1927 ( .in(\mat_kron/mult_40_G2/ab[4][0] ), .out(n1199) );
  oai22 U1928 ( .a(n1200), .b(n1199), .c(n2413), .d(n2414), .out(n1202) );
  aoi22 U1929 ( .a(n1202), .b(\mat_kron/mult_40_G2/ab[5][0] ), .c(n2415), .d(
        n1854), .out(n1207) );
  nand2 U1930 ( .a(\mat_kron/mult_40/ab[0][3] ), .b(
        \mat_kron/mult_40/ab[1][2] ), .out(n2416) );
  aoi22 U1931 ( .a(\mat_kron/mult_40/ab[2][2] ), .b(n1219), .c(n2417), .d(
        n1864), .out(n1222) );
  nand2 U1932 ( .a(\mat_kron/mult_40/ab[1][3] ), .b(
        \mat_kron/mult_40/ab[0][4] ), .out(n2418) );
  inv U1933 ( .in(\mat_kron/mult_40/ab[2][3] ), .out(n2419) );
  aoi22 U1934 ( .a(n2421), .b(\mat_kron/mult_40/ab[3][2] ), .c(n1220), .d(
        n1865), .out(n2420) );
  nand2 U1935 ( .a(\mat_kron/mult_40/ab[1][4] ), .b(
        \mat_kron/mult_40/ab[0][5] ), .out(n2422) );
  oai22 U1936 ( .a(n2418), .b(n2419), .c(n1212), .d(n1862), .out(n1217) );
  nand2 U1937 ( .a(\mat_kron/mult_40/ab[0][2] ), .b(
        \mat_kron/mult_40/ab[1][1] ), .out(n1229) );
  aoi22 U1938 ( .a(\mat_kron/mult_40/ab[2][1] ), .b(n2424), .c(n1227), .d(
        n1867), .out(n2423) );
  oai22 U1939 ( .a(n2423), .b(n2425), .c(n1230), .d(n1868), .out(n1233) );
  inv U1940 ( .in(\mat_kron/mult_40/ab[4][1] ), .out(n2426) );
  oai22 U1941 ( .a(n2427), .b(n2426), .c(n1232), .d(n1877), .out(n1235) );
  inv U1942 ( .in(\mat_kron/mult_40/ab[5][1] ), .out(n2428) );
  nand2 U1943 ( .a(\mat_kron/mult_40/ab[0][1] ), .b(
        \mat_kron/mult_40/ab[1][0] ), .out(n1238) );
  aoi22 U1944 ( .a(\mat_kron/mult_40/ab[2][0] ), .b(n2429), .c(n1236), .d(
        n1872), .out(n1241) );
  aoi22 U1945 ( .a(n2430), .b(\mat_kron/mult_40/ab[3][0] ), .c(n1239), .d(
        n1873), .out(n1244) );
  inv U1946 ( .in(\mat_kron/mult_40/ab[4][0] ), .out(n1243) );
  oai22 U1947 ( .a(n1244), .b(n1243), .c(n2431), .d(n2432), .out(n1246) );
  aoi22 U1948 ( .a(n1246), .b(\mat_kron/mult_40/ab[5][0] ), .c(n2433), .d(
        n1875), .out(n1251) );
  inv U1949 ( .in(A[9]), .out(n2434) );
  nor2 U1950 ( .a(A[8]), .b(\mat_sub/r102/B_AS [0]), .out(n191) );
  nor2 U1951 ( .a(A[0]), .b(\mat_sub/r106/B_AS [0]), .out(n195) );
  inv U1952 ( .in(A[1]), .out(n2435) );
  oai22 U1953 ( .a(n195), .b(n2436), .c(n1252), .d(n2435), .out(n1255) );
  aoi22 U1954 ( .a(n1255), .b(\mat_sub/r106/B_AS [2]), .c(n2437), .d(A[2]), 
        .out(n1258) );
  inv U1955 ( .in(A[3]), .out(n2438) );
  oai22 U1956 ( .a(n1258), .b(n1257), .c(n2439), .d(n2438), .out(n1260) );
  aoi22 U1957 ( .a(n1260), .b(\mat_sub/r106/B_AS [4]), .c(n2440), .d(A[4]), 
        .out(n1263) );
  inv U1958 ( .in(A[5]), .out(n2441) );
  oai22 U1959 ( .a(n1263), .b(n1262), .c(n2442), .d(n2441), .out(n1266) );
  nor2 U1960 ( .a(A[24]), .b(\mat_sub/r94/B_AS [0]), .out(n193) );
  inv U1961 ( .in(A[25]), .out(n2443) );
  oai22 U1962 ( .a(n193), .b(n2444), .c(n1267), .d(n2443), .out(n1270) );
  aoi22 U1963 ( .a(n1270), .b(\mat_sub/r94/B_AS [2]), .c(n2445), .d(A[26]), 
        .out(n1273) );
  inv U1964 ( .in(A[27]), .out(n2446) );
  oai22 U1965 ( .a(n1273), .b(n1272), .c(n2447), .d(n2446), .out(n1275) );
  aoi22 U1966 ( .a(n1275), .b(\mat_sub/r94/B_AS [4]), .c(n2448), .d(A[28]), 
        .out(n1278) );
  inv U1967 ( .in(A[29]), .out(n2449) );
  oai22 U1968 ( .a(n1278), .b(n1277), .c(n2450), .d(n2449), .out(n1281) );
  nor2 U1969 ( .a(A[16]), .b(\mat_sub/r98/B_AS [0]), .out(n189) );
  inv U1970 ( .in(A[17]), .out(n2451) );
  oai22 U1971 ( .a(n189), .b(n2452), .c(n1282), .d(n2451), .out(n1285) );
  aoi22 U1972 ( .a(n1285), .b(\mat_sub/r98/B_AS [2]), .c(n2453), .d(A[18]), 
        .out(n1288) );
  inv U1973 ( .in(A[19]), .out(n2454) );
  oai22 U1974 ( .a(n1288), .b(n1287), .c(n2455), .d(n2454), .out(n1290) );
  aoi22 U1975 ( .a(n1290), .b(\mat_sub/r98/B_AS [4]), .c(n2456), .d(A[20]), 
        .out(n1293) );
  inv U1976 ( .in(A[21]), .out(n2457) );
  oai22 U1977 ( .a(n1293), .b(n1292), .c(n2458), .d(n2457), .out(n1296) );
  aoi22 U1978 ( .a(n1298), .b(\mat_sub/r102/B_AS [1]), .c(n2459), .d(A[9]), 
        .out(n1301) );
  inv U1979 ( .in(\mat_sub/r102/B_AS [2]), .out(n1300) );
  aoi22 U1980 ( .a(n2460), .b(\mat_sub/r102/B_AS [2]), .c(n1299), .d(A[10]), 
        .out(n1304) );
  inv U1981 ( .in(A[11]), .out(n2461) );
  aoi22 U1982 ( .a(n2462), .b(\mat_sub/r102/B_AS [3]), .c(n1302), .d(A[11]), 
        .out(n1307) );
  inv U1983 ( .in(\mat_sub/r102/B_AS [4]), .out(n1306) );
  aoi22 U1984 ( .a(n2463), .b(\mat_sub/r102/B_AS [4]), .c(n1305), .d(A[12]), 
        .out(n1310) );
  inv U1985 ( .in(A[13]), .out(n2464) );
  inv U1986 ( .in(\mat_sub/r102/B_AS [5]), .out(n1309) );
  oai22 U1987 ( .a(n1310), .b(n1309), .c(n2465), .d(n2464), .out(n1313) );
  nand2 U1988 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[0] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[0] ), .out(n2466) );
  nand2 U1989 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[0] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[0] ), .out(n2467) );
  inv U1990 ( .in(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ), .out(n2468) );
  inv U1991 ( .in(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[3] ), .out(n2469) );
  inv U1992 ( .in(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ), .out(n2470) );
  inv U1993 ( .in(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[5] ), .out(n2471) );
  nand2 U1994 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[0] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[0] ), .out(n2472) );
  inv U1995 ( .in(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ), .out(n2473) );
  inv U1996 ( .in(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[3] ), .out(n2474) );
  inv U1997 ( .in(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ), .out(n2475) );
  inv U1998 ( .in(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[5] ), .out(n2476) );
  nand2 U1999 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[0] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[0] ), .out(n2477) );
  inv U2000 ( .in(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ), .out(n2478) );
  inv U2001 ( .in(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[3] ), .out(n2479) );
  inv U2002 ( .in(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ), .out(n2480) );
  inv U2003 ( .in(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[5] ), .out(n2481) );
  inv U2004 ( .in(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ), .out(n2482) );
  inv U2005 ( .in(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[3] ), .out(n2483) );
  inv U2006 ( .in(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ), .out(n2484) );
  inv U2007 ( .in(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[5] ), .out(n2485) );
  nand2 U2008 ( .a(\mat_add/r102/B_AS [0]), .b(A[8]), .out(n2486) );
  inv U2009 ( .in(\mat_add/r102/B_AS [1]), .out(n2487) );
  nand2 U2010 ( .a(\mat_add/r106/B_AS [0]), .b(A[0]), .out(n2488) );
  inv U2011 ( .in(\mat_add/r106/B_AS [1]), .out(n2489) );
  inv U2012 ( .in(\mat_add/r106/B_AS [3]), .out(n2490) );
  inv U2013 ( .in(\mat_add/r106/B_AS [5]), .out(n2491) );
  nand2 U2014 ( .a(\mat_add/r94/B_AS [0]), .b(A[24]), .out(n2492) );
  inv U2015 ( .in(\mat_add/r94/B_AS [1]), .out(n2493) );
  inv U2016 ( .in(\mat_add/r94/B_AS [3]), .out(n2494) );
  inv U2017 ( .in(\mat_add/r94/B_AS [5]), .out(n2495) );
  nand2 U2018 ( .a(\mat_add/r98/B_AS [0]), .b(A[16]), .out(n2496) );
  inv U2019 ( .in(\mat_add/r98/B_AS [1]), .out(n2497) );
  inv U2020 ( .in(\mat_add/r98/B_AS [3]), .out(n2498) );
  inv U2021 ( .in(\mat_add/r98/B_AS [5]), .out(n2499) );
  inv U2022 ( .in(\mat_add/r102/B_AS [3]), .out(n2500) );
  inv U2023 ( .in(\mat_add/r102/B_AS [5]), .out(n2501) );
  xor2 U2024 ( .a(n2503), .b(n2504), .out(n2502) );
  xor2 U2025 ( .a(n236), .b(n2505), .out(\mat_mul/mult_37_G2_G2_G2/A1[4] ) );
  xor2 U2026 ( .a(n2018), .b(n2506), .out(\mat_mul/mult_37_G2_G2_G2/A1[2] ) );
  xor2 U2027 ( .a(n1389), .b(n2507), .out(\mat_mul/mult_37_G2_G2_G2/A1[0] ) );
  xor2 U2028 ( .a(n2509), .b(n2510), .out(n2508) );
  xor2 U2029 ( .a(n280), .b(n2511), .out(\mat_mul/mult_37_G2_G2_G1/A1[4] ) );
  xor2 U2030 ( .a(n2036), .b(n2512), .out(\mat_mul/mult_37_G2_G2_G1/A1[2] ) );
  xor2 U2031 ( .a(n1410), .b(n2513), .out(\mat_mul/mult_37_G2_G2_G1/A1[0] ) );
  xor2 U2032 ( .a(n2515), .b(n2516), .out(n2514) );
  xor2 U2033 ( .a(n324), .b(n2517), .out(\mat_mul/mult_37_G2_G2/A1[4] ) );
  xor2 U2034 ( .a(n2054), .b(n2518), .out(\mat_mul/mult_37_G2_G2/A1[2] ) );
  xor2 U2035 ( .a(n1431), .b(n2519), .out(\mat_mul/mult_37_G2_G2/A1[0] ) );
  xor2 U2036 ( .a(n2521), .b(n2522), .out(n2520) );
  xor2 U2037 ( .a(n368), .b(n2523), .out(\mat_mul/mult_37_G2_G1_G2/A1[4] ) );
  xor2 U2038 ( .a(n2072), .b(n2524), .out(\mat_mul/mult_37_G2_G1_G2/A1[2] ) );
  xor2 U2039 ( .a(n1452), .b(n2525), .out(\mat_mul/mult_37_G2_G1_G2/A1[0] ) );
  xor2 U2040 ( .a(n2527), .b(n2528), .out(n2526) );
  xor2 U2041 ( .a(n412), .b(n2529), .out(\mat_mul/mult_37_G2_G1_G1/A1[4] ) );
  xor2 U2042 ( .a(n2090), .b(n2530), .out(\mat_mul/mult_37_G2_G1_G1/A1[2] ) );
  xor2 U2043 ( .a(n1473), .b(n2531), .out(\mat_mul/mult_37_G2_G1_G1/A1[0] ) );
  xor2 U2044 ( .a(n2533), .b(n2534), .out(n2532) );
  xor2 U2045 ( .a(n456), .b(n2535), .out(\mat_mul/mult_37_G2_G1/A1[4] ) );
  xor2 U2046 ( .a(n2108), .b(n2536), .out(\mat_mul/mult_37_G2_G1/A1[2] ) );
  xor2 U2047 ( .a(n1494), .b(n2537), .out(\mat_mul/mult_37_G2_G1/A1[0] ) );
  xor2 U2048 ( .a(n2539), .b(n2540), .out(n2538) );
  xor2 U2049 ( .a(n500), .b(n2541), .out(\mat_mul/mult_37_G2/A1[4] ) );
  xor2 U2050 ( .a(n2126), .b(n2542), .out(\mat_mul/mult_37_G2/A1[2] ) );
  xor2 U2051 ( .a(n1515), .b(n2543), .out(\mat_mul/mult_37_G2/A1[0] ) );
  xor2 U2052 ( .a(n2545), .b(n2546), .out(n2544) );
  xor2 U2053 ( .a(n544), .b(n2547), .out(\mat_mul/mult_37/A1[4] ) );
  xor2 U2054 ( .a(n2144), .b(n2548), .out(\mat_mul/mult_37/A1[2] ) );
  xor2 U2055 ( .a(n1536), .b(n2549), .out(\mat_mul/mult_37/A1[0] ) );
  xor2 U2056 ( .a(n2551), .b(n2552), .out(n2550) );
  xor2 U2057 ( .a(n588), .b(n2553), .out(\mat_kron/mult_40_G2_G2_G2_G2/A1[4] )
         );
  xor2 U2058 ( .a(n2162), .b(n2554), .out(\mat_kron/mult_40_G2_G2_G2_G2/A1[2] ) );
  xor2 U2059 ( .a(n1557), .b(n2555), .out(\mat_kron/mult_40_G2_G2_G2_G2/A1[0] ) );
  xor2 U2060 ( .a(n2557), .b(n2558), .out(n2556) );
  xor2 U2061 ( .a(n632), .b(n2559), .out(\mat_kron/mult_40_G2_G2_G2_G1/A1[4] )
         );
  xor2 U2062 ( .a(n2180), .b(n2560), .out(\mat_kron/mult_40_G2_G2_G2_G1/A1[2] ) );
  xor2 U2063 ( .a(n1578), .b(n2561), .out(\mat_kron/mult_40_G2_G2_G2_G1/A1[0] ) );
  xor2 U2064 ( .a(n2563), .b(n2564), .out(n2562) );
  xor2 U2065 ( .a(n676), .b(n2565), .out(\mat_kron/mult_40_G2_G2_G2/A1[4] ) );
  xor2 U2066 ( .a(n2198), .b(n2566), .out(\mat_kron/mult_40_G2_G2_G2/A1[2] )
         );
  xor2 U2067 ( .a(n1599), .b(n2567), .out(\mat_kron/mult_40_G2_G2_G2/A1[0] )
         );
  xor2 U2068 ( .a(n2569), .b(n2570), .out(n2568) );
  xor2 U2069 ( .a(n720), .b(n2571), .out(\mat_kron/mult_40_G2_G2_G1_G2/A1[4] )
         );
  xor2 U2070 ( .a(n2216), .b(n2572), .out(\mat_kron/mult_40_G2_G2_G1_G2/A1[2] ) );
  xor2 U2071 ( .a(n1620), .b(n2573), .out(\mat_kron/mult_40_G2_G2_G1_G2/A1[0] ) );
  xor2 U2072 ( .a(n2575), .b(n2576), .out(n2574) );
  xor2 U2073 ( .a(n764), .b(n2577), .out(\mat_kron/mult_40_G2_G2_G1_G1/A1[4] )
         );
  xor2 U2074 ( .a(n2234), .b(n2578), .out(\mat_kron/mult_40_G2_G2_G1_G1/A1[2] ) );
  xor2 U2075 ( .a(n1641), .b(n2579), .out(\mat_kron/mult_40_G2_G2_G1_G1/A1[0] ) );
  xor2 U2076 ( .a(n2581), .b(n2582), .out(n2580) );
  xor2 U2077 ( .a(n808), .b(n2583), .out(\mat_kron/mult_40_G2_G2_G1/A1[4] ) );
  xor2 U2078 ( .a(n2252), .b(n2584), .out(\mat_kron/mult_40_G2_G2_G1/A1[2] )
         );
  xor2 U2079 ( .a(n1662), .b(n2585), .out(\mat_kron/mult_40_G2_G2_G1/A1[0] )
         );
  xor2 U2080 ( .a(n2587), .b(n2588), .out(n2586) );
  xor2 U2081 ( .a(n852), .b(n2589), .out(\mat_kron/mult_40_G2_G2/A1[4] ) );
  xor2 U2082 ( .a(n2270), .b(n2590), .out(\mat_kron/mult_40_G2_G2/A1[2] ) );
  xor2 U2083 ( .a(n1683), .b(n2591), .out(\mat_kron/mult_40_G2_G2/A1[0] ) );
  xor2 U2084 ( .a(n2593), .b(n2594), .out(n2592) );
  xor2 U2085 ( .a(n896), .b(n2595), .out(\mat_kron/mult_40_G2_G1_G2_G2/A1[4] )
         );
  xor2 U2086 ( .a(n2288), .b(n2596), .out(\mat_kron/mult_40_G2_G1_G2_G2/A1[2] ) );
  xor2 U2087 ( .a(n1704), .b(n2597), .out(\mat_kron/mult_40_G2_G1_G2_G2/A1[0] ) );
  xor2 U2088 ( .a(n2599), .b(n2600), .out(n2598) );
  xor2 U2089 ( .a(n940), .b(n2601), .out(\mat_kron/mult_40_G2_G1_G2_G1/A1[4] )
         );
  xor2 U2090 ( .a(n2306), .b(n2602), .out(\mat_kron/mult_40_G2_G1_G2_G1/A1[2] ) );
  xor2 U2091 ( .a(n1725), .b(n2603), .out(\mat_kron/mult_40_G2_G1_G2_G1/A1[0] ) );
  xor2 U2092 ( .a(n2605), .b(n2606), .out(n2604) );
  xor2 U2093 ( .a(n984), .b(n2607), .out(\mat_kron/mult_40_G2_G1_G2/A1[4] ) );
  xor2 U2094 ( .a(n2324), .b(n2608), .out(\mat_kron/mult_40_G2_G1_G2/A1[2] )
         );
  xor2 U2095 ( .a(n1746), .b(n2609), .out(\mat_kron/mult_40_G2_G1_G2/A1[0] )
         );
  xor2 U2096 ( .a(n2611), .b(n2612), .out(n2610) );
  xor2 U2097 ( .a(n1028), .b(n2613), .out(\mat_kron/mult_40_G2_G1_G1_G2/A1[4] ) );
  xor2 U2098 ( .a(n2342), .b(n2614), .out(\mat_kron/mult_40_G2_G1_G1_G2/A1[2] ) );
  xor2 U2099 ( .a(n1767), .b(n2615), .out(\mat_kron/mult_40_G2_G1_G1_G2/A1[0] ) );
  xor2 U2100 ( .a(n2617), .b(n2618), .out(n2616) );
  xor2 U2101 ( .a(n1072), .b(n2619), .out(\mat_kron/mult_40_G2_G1_G1_G1/A1[4] ) );
  xor2 U2102 ( .a(n2360), .b(n2620), .out(\mat_kron/mult_40_G2_G1_G1_G1/A1[2] ) );
  xor2 U2103 ( .a(n1788), .b(n2621), .out(\mat_kron/mult_40_G2_G1_G1_G1/A1[0] ) );
  xor2 U2104 ( .a(n2623), .b(n2624), .out(n2622) );
  xor2 U2105 ( .a(n1116), .b(n2625), .out(\mat_kron/mult_40_G2_G1_G1/A1[4] )
         );
  xor2 U2106 ( .a(n2378), .b(n2626), .out(\mat_kron/mult_40_G2_G1_G1/A1[2] )
         );
  xor2 U2107 ( .a(n1809), .b(n2627), .out(\mat_kron/mult_40_G2_G1_G1/A1[0] )
         );
  xor2 U2108 ( .a(n2629), .b(n2630), .out(n2628) );
  xor2 U2109 ( .a(n1160), .b(n2631), .out(\mat_kron/mult_40_G2_G1/A1[4] ) );
  xor2 U2110 ( .a(n2396), .b(n2632), .out(\mat_kron/mult_40_G2_G1/A1[2] ) );
  xor2 U2111 ( .a(n1830), .b(n2633), .out(\mat_kron/mult_40_G2_G1/A1[0] ) );
  xor2 U2112 ( .a(n2635), .b(n2636), .out(n2634) );
  xor2 U2113 ( .a(n1204), .b(n2637), .out(\mat_kron/mult_40_G2/A1[4] ) );
  xor2 U2114 ( .a(n2414), .b(n2638), .out(\mat_kron/mult_40_G2/A1[2] ) );
  xor2 U2115 ( .a(n1851), .b(n2639), .out(\mat_kron/mult_40_G2/A1[0] ) );
  xor2 U2116 ( .a(n2641), .b(n2642), .out(n2640) );
  xor2 U2117 ( .a(n1248), .b(n2643), .out(\mat_kron/mult_40/A1[4] ) );
  xor2 U2118 ( .a(n2432), .b(n2644), .out(\mat_kron/mult_40/A1[2] ) );
  xor2 U2119 ( .a(n1872), .b(n2645), .out(\mat_kron/mult_40/A1[0] ) );
  xor2 U2120 ( .a(n1339), .b(n2646), .out(m_mul[9]) );
  xor2 U2121 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[0] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[0] ), .out(m_mul[8]) );
  xor2 U2122 ( .a(n1324), .b(n2647), .out(m_mul[25]) );
  xor2 U2123 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[0] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[0] ), .out(m_mul[24]) );
  xor2 U2124 ( .a(n1316), .b(n2648), .out(m_mul[1]) );
  xor2 U2125 ( .a(n1332), .b(n2649), .out(m_mul[17]) );
  xor2 U2126 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[0] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[0] ), .out(m_mul[16]) );
  xor2 U2127 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[0] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[0] ), .out(m_mul[0]) );
  xor2 U2128 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G2_G2/ab[1][0] ), .out(m_kro[9]) );
  xor2 U2129 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[1][0] ), .out(m_kro[97]) );
  xor2 U2130 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G1_G1/ab[1][0] ), .out(m_kro[89]) );
  xor2 U2131 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[1][0] ), .out(m_kro[81]) );
  xor2 U2132 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G2_G1/ab[1][0] ), .out(m_kro[73]) );
  xor2 U2133 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[1][0] ), .out(m_kro[65]) );
  xor2 U2134 ( .a(\mat_kron/mult_40_G2/ab[0][1] ), .b(
        \mat_kron/mult_40_G2/ab[1][0] ), .out(m_kro[57]) );
  xor2 U2135 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[1][0] ), .out(m_kro[49]) );
  xor2 U2136 ( .a(\mat_kron/mult_40_G2_G2/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G2/ab[1][0] ), .out(m_kro[41]) );
  xor2 U2137 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[1][0] ), .out(m_kro[33]) );
  xor2 U2138 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G1_G2/ab[1][0] ), .out(m_kro[25]) );
  xor2 U2139 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[1][0] ), .out(m_kro[1]) );
  xor2 U2140 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[1][0] ), .out(m_kro[17]) );
  xor2 U2141 ( .a(\mat_kron/mult_40/ab[0][1] ), .b(\mat_kron/mult_40/ab[1][0] ), .out(m_kro[121]) );
  xor2 U2142 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[1][0] ), .out(m_kro[113]) );
  xor2 U2143 ( .a(\mat_kron/mult_40_G2_G1/ab[0][1] ), .b(
        \mat_kron/mult_40_G2_G1/ab[1][0] ), .out(m_kro[105]) );
  xor2 U2144 ( .a(n2487), .b(n2650), .out(m_add[9]) );
  xor2 U2145 ( .a(A[8]), .b(\mat_add/r102/B_AS [0]), .out(m_add[8]) );
  xor2 U2146 ( .a(n2493), .b(n2651), .out(m_add[25]) );
  xor2 U2147 ( .a(A[24]), .b(\mat_add/r94/B_AS [0]), .out(m_add[24]) );
  xor2 U2148 ( .a(n2489), .b(n2652), .out(m_add[1]) );
  xor2 U2149 ( .a(n2497), .b(n2653), .out(m_add[17]) );
  xor2 U2150 ( .a(A[16]), .b(\mat_add/r98/B_AS [0]), .out(m_add[16]) );
  xor2 U2151 ( .a(A[0]), .b(\mat_add/r106/B_AS [0]), .out(m_add[0]) );
  xor2 U2152 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[0][7] ), .b(
        \mat_mul/mult_37_G2_G2_G2/ab[1][6] ), .out(n2654) );
  xor2 U2153 ( .a(n164), .b(\mat_mul/mult_37_G2_G2_G2/ab[2][5] ), .out(n2655)
         );
  xor2 U2154 ( .a(n2654), .b(n2655), .out(n2503) );
  xor2 U2155 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[3][4] ), .b(
        \mat_mul/mult_37_G2_G2_G2/ab[4][3] ), .out(n2656) );
  xor2 U2156 ( .a(n196), .b(n202), .out(n2657) );
  xor2 U2157 ( .a(n2656), .b(n2657), .out(n2504) );
  xor2 U2158 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[5][2] ), .b(
        \mat_mul/mult_37_G2_G2_G2/ab[6][1] ), .out(n2658) );
  xor2 U2159 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[7][0] ), .b(n211), .out(n2659)
         );
  xor2 U2160 ( .a(n2658), .b(n2659), .out(n1396) );
  xor2 U2161 ( .a(n238), .b(n2660), .out(n2505) );
  xor2 U2162 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[4][0] ), .b(n232), .out(n2506)
         );
  xor2 U2163 ( .a(n2015), .b(\mat_mul/mult_37_G2_G2_G2/ab[2][0] ), .out(n2507)
         );
  xor2 U2164 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[0][7] ), .b(
        \mat_mul/mult_37_G2_G2_G1/ab[1][6] ), .out(n2661) );
  xor2 U2165 ( .a(n168), .b(\mat_mul/mult_37_G2_G2_G1/ab[2][5] ), .out(n2662)
         );
  xor2 U2166 ( .a(n2661), .b(n2662), .out(n2509) );
  xor2 U2167 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[3][4] ), .b(
        \mat_mul/mult_37_G2_G2_G1/ab[4][3] ), .out(n2663) );
  xor2 U2168 ( .a(n240), .b(n246), .out(n2664) );
  xor2 U2169 ( .a(n2663), .b(n2664), .out(n2510) );
  xor2 U2170 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[5][2] ), .b(
        \mat_mul/mult_37_G2_G2_G1/ab[6][1] ), .out(n2665) );
  xor2 U2171 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[7][0] ), .b(n255), .out(n2666)
         );
  xor2 U2172 ( .a(n2665), .b(n2666), .out(n1417) );
  xor2 U2173 ( .a(n282), .b(n2667), .out(n2511) );
  xor2 U2174 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[4][0] ), .b(n276), .out(n2512)
         );
  xor2 U2175 ( .a(n2033), .b(\mat_mul/mult_37_G2_G2_G1/ab[2][0] ), .out(n2513)
         );
  xor2 U2176 ( .a(\mat_mul/mult_37_G2_G2/ab[0][7] ), .b(
        \mat_mul/mult_37_G2_G2/ab[1][6] ), .out(n2668) );
  xor2 U2177 ( .a(n165), .b(\mat_mul/mult_37_G2_G2/ab[2][5] ), .out(n2669) );
  xor2 U2178 ( .a(n2668), .b(n2669), .out(n2515) );
  xor2 U2179 ( .a(\mat_mul/mult_37_G2_G2/ab[3][4] ), .b(
        \mat_mul/mult_37_G2_G2/ab[4][3] ), .out(n2670) );
  xor2 U2180 ( .a(n284), .b(n290), .out(n2671) );
  xor2 U2181 ( .a(n2670), .b(n2671), .out(n2516) );
  xor2 U2182 ( .a(\mat_mul/mult_37_G2_G2/ab[5][2] ), .b(
        \mat_mul/mult_37_G2_G2/ab[6][1] ), .out(n2672) );
  xor2 U2183 ( .a(\mat_mul/mult_37_G2_G2/ab[7][0] ), .b(n299), .out(n2673) );
  xor2 U2184 ( .a(n2672), .b(n2673), .out(n1438) );
  xor2 U2185 ( .a(n326), .b(n2674), .out(n2517) );
  xor2 U2186 ( .a(\mat_mul/mult_37_G2_G2/ab[4][0] ), .b(n320), .out(n2518) );
  xor2 U2187 ( .a(n2051), .b(\mat_mul/mult_37_G2_G2/ab[2][0] ), .out(n2519) );
  xor2 U2188 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[0][7] ), .b(
        \mat_mul/mult_37_G2_G1_G2/ab[1][6] ), .out(n2675) );
  xor2 U2189 ( .a(n166), .b(\mat_mul/mult_37_G2_G1_G2/ab[2][5] ), .out(n2676)
         );
  xor2 U2190 ( .a(n2675), .b(n2676), .out(n2521) );
  xor2 U2191 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[3][4] ), .b(
        \mat_mul/mult_37_G2_G1_G2/ab[4][3] ), .out(n2677) );
  xor2 U2192 ( .a(n328), .b(n334), .out(n2678) );
  xor2 U2193 ( .a(n2677), .b(n2678), .out(n2522) );
  xor2 U2194 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[5][2] ), .b(
        \mat_mul/mult_37_G2_G1_G2/ab[6][1] ), .out(n2679) );
  xor2 U2195 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[7][0] ), .b(n343), .out(n2680)
         );
  xor2 U2196 ( .a(n2679), .b(n2680), .out(n1459) );
  xor2 U2197 ( .a(n370), .b(n2681), .out(n2523) );
  xor2 U2198 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[4][0] ), .b(n364), .out(n2524)
         );
  xor2 U2199 ( .a(n2069), .b(\mat_mul/mult_37_G2_G1_G2/ab[2][0] ), .out(n2525)
         );
  xor2 U2200 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[0][7] ), .b(
        \mat_mul/mult_37_G2_G1_G1/ab[1][6] ), .out(n2682) );
  xor2 U2201 ( .a(n170), .b(\mat_mul/mult_37_G2_G1_G1/ab[2][5] ), .out(n2683)
         );
  xor2 U2202 ( .a(n2682), .b(n2683), .out(n2527) );
  xor2 U2203 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[3][4] ), .b(
        \mat_mul/mult_37_G2_G1_G1/ab[4][3] ), .out(n2684) );
  xor2 U2204 ( .a(n372), .b(n378), .out(n2685) );
  xor2 U2205 ( .a(n2684), .b(n2685), .out(n2528) );
  xor2 U2206 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[5][2] ), .b(
        \mat_mul/mult_37_G2_G1_G1/ab[6][1] ), .out(n2686) );
  xor2 U2207 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[7][0] ), .b(n387), .out(n2687)
         );
  xor2 U2208 ( .a(n2686), .b(n2687), .out(n1480) );
  xor2 U2209 ( .a(n414), .b(n2688), .out(n2529) );
  xor2 U2210 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[4][0] ), .b(n408), .out(n2530)
         );
  xor2 U2211 ( .a(n2087), .b(\mat_mul/mult_37_G2_G1_G1/ab[2][0] ), .out(n2531)
         );
  xor2 U2212 ( .a(\mat_mul/mult_37_G2_G1/ab[0][7] ), .b(
        \mat_mul/mult_37_G2_G1/ab[1][6] ), .out(n2689) );
  xor2 U2213 ( .a(n169), .b(\mat_mul/mult_37_G2_G1/ab[2][5] ), .out(n2690) );
  xor2 U2214 ( .a(n2689), .b(n2690), .out(n2533) );
  xor2 U2215 ( .a(\mat_mul/mult_37_G2_G1/ab[3][4] ), .b(
        \mat_mul/mult_37_G2_G1/ab[4][3] ), .out(n2691) );
  xor2 U2216 ( .a(n416), .b(n422), .out(n2692) );
  xor2 U2217 ( .a(n2691), .b(n2692), .out(n2534) );
  xor2 U2218 ( .a(\mat_mul/mult_37_G2_G1/ab[5][2] ), .b(
        \mat_mul/mult_37_G2_G1/ab[6][1] ), .out(n2693) );
  xor2 U2219 ( .a(\mat_mul/mult_37_G2_G1/ab[7][0] ), .b(n431), .out(n2694) );
  xor2 U2220 ( .a(n2693), .b(n2694), .out(n1501) );
  xor2 U2221 ( .a(n458), .b(n2695), .out(n2535) );
  xor2 U2222 ( .a(\mat_mul/mult_37_G2_G1/ab[4][0] ), .b(n452), .out(n2536) );
  xor2 U2223 ( .a(n2105), .b(\mat_mul/mult_37_G2_G1/ab[2][0] ), .out(n2537) );
  xor2 U2224 ( .a(\mat_mul/mult_37_G2/ab[0][7] ), .b(
        \mat_mul/mult_37_G2/ab[1][6] ), .out(n2696) );
  xor2 U2225 ( .a(n167), .b(\mat_mul/mult_37_G2/ab[2][5] ), .out(n2697) );
  xor2 U2226 ( .a(n2696), .b(n2697), .out(n2539) );
  xor2 U2227 ( .a(\mat_mul/mult_37_G2/ab[3][4] ), .b(
        \mat_mul/mult_37_G2/ab[4][3] ), .out(n2698) );
  xor2 U2228 ( .a(n460), .b(n466), .out(n2699) );
  xor2 U2229 ( .a(n2698), .b(n2699), .out(n2540) );
  xor2 U2230 ( .a(\mat_mul/mult_37_G2/ab[5][2] ), .b(
        \mat_mul/mult_37_G2/ab[6][1] ), .out(n2700) );
  xor2 U2231 ( .a(\mat_mul/mult_37_G2/ab[7][0] ), .b(n475), .out(n2701) );
  xor2 U2232 ( .a(n2700), .b(n2701), .out(n1522) );
  xor2 U2233 ( .a(n502), .b(n2702), .out(n2541) );
  xor2 U2234 ( .a(\mat_mul/mult_37_G2/ab[4][0] ), .b(n496), .out(n2542) );
  xor2 U2235 ( .a(n2123), .b(\mat_mul/mult_37_G2/ab[2][0] ), .out(n2543) );
  xor2 U2236 ( .a(\mat_mul/mult_37/ab[0][7] ), .b(\mat_mul/mult_37/ab[1][6] ), 
        .out(n2703) );
  xor2 U2237 ( .a(n171), .b(\mat_mul/mult_37/ab[2][5] ), .out(n2704) );
  xor2 U2238 ( .a(n2703), .b(n2704), .out(n2545) );
  xor2 U2239 ( .a(\mat_mul/mult_37/ab[3][4] ), .b(\mat_mul/mult_37/ab[4][3] ), 
        .out(n2705) );
  xor2 U2240 ( .a(n504), .b(n510), .out(n2706) );
  xor2 U2241 ( .a(n2705), .b(n2706), .out(n2546) );
  xor2 U2242 ( .a(\mat_mul/mult_37/ab[5][2] ), .b(\mat_mul/mult_37/ab[6][1] ), 
        .out(n2707) );
  xor2 U2243 ( .a(\mat_mul/mult_37/ab[7][0] ), .b(n519), .out(n2708) );
  xor2 U2244 ( .a(n2707), .b(n2708), .out(n1543) );
  xor2 U2245 ( .a(n546), .b(n2709), .out(n2547) );
  xor2 U2246 ( .a(\mat_mul/mult_37/ab[4][0] ), .b(n540), .out(n2548) );
  xor2 U2247 ( .a(n2141), .b(\mat_mul/mult_37/ab[2][0] ), .out(n2549) );
  xor2 U2248 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[0][7] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[1][6] ), .out(n2710) );
  xor2 U2249 ( .a(n172), .b(\mat_kron/mult_40_G2_G2_G2_G2/ab[2][5] ), .out(
        n2711) );
  xor2 U2250 ( .a(n2710), .b(n2711), .out(n2551) );
  xor2 U2251 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[3][4] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[4][3] ), .out(n2712) );
  xor2 U2252 ( .a(n548), .b(n554), .out(n2713) );
  xor2 U2253 ( .a(n2712), .b(n2713), .out(n2552) );
  xor2 U2254 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[5][2] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G2/ab[6][1] ), .out(n2714) );
  xor2 U2255 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[7][0] ), .b(n563), .out(
        n2715) );
  xor2 U2256 ( .a(n2714), .b(n2715), .out(n1564) );
  xor2 U2257 ( .a(n590), .b(n2716), .out(n2553) );
  xor2 U2258 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[4][0] ), .b(n584), .out(
        n2554) );
  xor2 U2259 ( .a(n2159), .b(\mat_kron/mult_40_G2_G2_G2_G2/ab[2][0] ), .out(
        n2555) );
  xor2 U2260 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[0][7] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[1][6] ), .out(n2717) );
  xor2 U2261 ( .a(n180), .b(\mat_kron/mult_40_G2_G2_G2_G1/ab[2][5] ), .out(
        n2718) );
  xor2 U2262 ( .a(n2717), .b(n2718), .out(n2557) );
  xor2 U2263 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[3][4] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[4][3] ), .out(n2719) );
  xor2 U2264 ( .a(n592), .b(n598), .out(n2720) );
  xor2 U2265 ( .a(n2719), .b(n2720), .out(n2558) );
  xor2 U2266 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[5][2] ), .b(
        \mat_kron/mult_40_G2_G2_G2_G1/ab[6][1] ), .out(n2721) );
  xor2 U2267 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[7][0] ), .b(n607), .out(
        n2722) );
  xor2 U2268 ( .a(n2721), .b(n2722), .out(n1585) );
  xor2 U2269 ( .a(n634), .b(n2723), .out(n2559) );
  xor2 U2270 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[4][0] ), .b(n628), .out(
        n2560) );
  xor2 U2271 ( .a(n2177), .b(\mat_kron/mult_40_G2_G2_G2_G1/ab[2][0] ), .out(
        n2561) );
  xor2 U2272 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[0][7] ), .b(
        \mat_kron/mult_40_G2_G2_G2/ab[1][6] ), .out(n2724) );
  xor2 U2273 ( .a(n173), .b(\mat_kron/mult_40_G2_G2_G2/ab[2][5] ), .out(n2725)
         );
  xor2 U2274 ( .a(n2724), .b(n2725), .out(n2563) );
  xor2 U2275 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[3][4] ), .b(
        \mat_kron/mult_40_G2_G2_G2/ab[4][3] ), .out(n2726) );
  xor2 U2276 ( .a(n636), .b(n642), .out(n2727) );
  xor2 U2277 ( .a(n2726), .b(n2727), .out(n2564) );
  xor2 U2278 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[5][2] ), .b(
        \mat_kron/mult_40_G2_G2_G2/ab[6][1] ), .out(n2728) );
  xor2 U2279 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[7][0] ), .b(n651), .out(n2729)
         );
  xor2 U2280 ( .a(n2728), .b(n2729), .out(n1606) );
  xor2 U2281 ( .a(n678), .b(n2730), .out(n2565) );
  xor2 U2282 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[4][0] ), .b(n672), .out(n2566)
         );
  xor2 U2283 ( .a(n2195), .b(\mat_kron/mult_40_G2_G2_G2/ab[2][0] ), .out(n2567) );
  xor2 U2284 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[0][7] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[1][6] ), .out(n2731) );
  xor2 U2285 ( .a(n176), .b(\mat_kron/mult_40_G2_G2_G1_G2/ab[2][5] ), .out(
        n2732) );
  xor2 U2286 ( .a(n2731), .b(n2732), .out(n2569) );
  xor2 U2287 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[3][4] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[4][3] ), .out(n2733) );
  xor2 U2288 ( .a(n680), .b(n686), .out(n2734) );
  xor2 U2289 ( .a(n2733), .b(n2734), .out(n2570) );
  xor2 U2290 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[5][2] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G2/ab[6][1] ), .out(n2735) );
  xor2 U2291 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[7][0] ), .b(n695), .out(
        n2736) );
  xor2 U2292 ( .a(n2735), .b(n2736), .out(n1627) );
  xor2 U2293 ( .a(n722), .b(n2737), .out(n2571) );
  xor2 U2294 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[4][0] ), .b(n716), .out(
        n2572) );
  xor2 U2295 ( .a(n2213), .b(\mat_kron/mult_40_G2_G2_G1_G2/ab[2][0] ), .out(
        n2573) );
  xor2 U2296 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[0][7] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[1][6] ), .out(n2738) );
  xor2 U2297 ( .a(n184), .b(\mat_kron/mult_40_G2_G2_G1_G1/ab[2][5] ), .out(
        n2739) );
  xor2 U2298 ( .a(n2738), .b(n2739), .out(n2575) );
  xor2 U2299 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[3][4] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[4][3] ), .out(n2740) );
  xor2 U2300 ( .a(n724), .b(n730), .out(n2741) );
  xor2 U2301 ( .a(n2740), .b(n2741), .out(n2576) );
  xor2 U2302 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[5][2] ), .b(
        \mat_kron/mult_40_G2_G2_G1_G1/ab[6][1] ), .out(n2742) );
  xor2 U2303 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[7][0] ), .b(n739), .out(
        n2743) );
  xor2 U2304 ( .a(n2742), .b(n2743), .out(n1648) );
  xor2 U2305 ( .a(n766), .b(n2744), .out(n2577) );
  xor2 U2306 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[4][0] ), .b(n760), .out(
        n2578) );
  xor2 U2307 ( .a(n2231), .b(\mat_kron/mult_40_G2_G2_G1_G1/ab[2][0] ), .out(
        n2579) );
  xor2 U2308 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[0][7] ), .b(
        \mat_kron/mult_40_G2_G2_G1/ab[1][6] ), .out(n2745) );
  xor2 U2309 ( .a(n181), .b(\mat_kron/mult_40_G2_G2_G1/ab[2][5] ), .out(n2746)
         );
  xor2 U2310 ( .a(n2745), .b(n2746), .out(n2581) );
  xor2 U2311 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[3][4] ), .b(
        \mat_kron/mult_40_G2_G2_G1/ab[4][3] ), .out(n2747) );
  xor2 U2312 ( .a(n768), .b(n774), .out(n2748) );
  xor2 U2313 ( .a(n2747), .b(n2748), .out(n2582) );
  xor2 U2314 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[5][2] ), .b(
        \mat_kron/mult_40_G2_G2_G1/ab[6][1] ), .out(n2749) );
  xor2 U2315 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[7][0] ), .b(n783), .out(n2750)
         );
  xor2 U2316 ( .a(n2749), .b(n2750), .out(n1669) );
  xor2 U2317 ( .a(n810), .b(n2751), .out(n2583) );
  xor2 U2318 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[4][0] ), .b(n804), .out(n2584)
         );
  xor2 U2319 ( .a(n2249), .b(\mat_kron/mult_40_G2_G2_G1/ab[2][0] ), .out(n2585) );
  xor2 U2320 ( .a(\mat_kron/mult_40_G2_G2/ab[0][7] ), .b(
        \mat_kron/mult_40_G2_G2/ab[1][6] ), .out(n2752) );
  xor2 U2321 ( .a(n175), .b(\mat_kron/mult_40_G2_G2/ab[2][5] ), .out(n2753) );
  xor2 U2322 ( .a(n2752), .b(n2753), .out(n2587) );
  xor2 U2323 ( .a(\mat_kron/mult_40_G2_G2/ab[3][4] ), .b(
        \mat_kron/mult_40_G2_G2/ab[4][3] ), .out(n2754) );
  xor2 U2324 ( .a(n812), .b(n818), .out(n2755) );
  xor2 U2325 ( .a(n2754), .b(n2755), .out(n2588) );
  xor2 U2326 ( .a(\mat_kron/mult_40_G2_G2/ab[5][2] ), .b(
        \mat_kron/mult_40_G2_G2/ab[6][1] ), .out(n2756) );
  xor2 U2327 ( .a(\mat_kron/mult_40_G2_G2/ab[7][0] ), .b(n827), .out(n2757) );
  xor2 U2328 ( .a(n2756), .b(n2757), .out(n1690) );
  xor2 U2329 ( .a(n854), .b(n2758), .out(n2589) );
  xor2 U2330 ( .a(\mat_kron/mult_40_G2_G2/ab[4][0] ), .b(n848), .out(n2590) );
  xor2 U2331 ( .a(n2267), .b(\mat_kron/mult_40_G2_G2/ab[2][0] ), .out(n2591)
         );
  xor2 U2332 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[0][7] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[1][6] ), .out(n2759) );
  xor2 U2333 ( .a(n174), .b(\mat_kron/mult_40_G2_G1_G2_G2/ab[2][5] ), .out(
        n2760) );
  xor2 U2334 ( .a(n2759), .b(n2760), .out(n2593) );
  xor2 U2335 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[3][4] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[4][3] ), .out(n2761) );
  xor2 U2336 ( .a(n856), .b(n862), .out(n2762) );
  xor2 U2337 ( .a(n2761), .b(n2762), .out(n2594) );
  xor2 U2338 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[5][2] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G2/ab[6][1] ), .out(n2763) );
  xor2 U2339 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[7][0] ), .b(n871), .out(
        n2764) );
  xor2 U2340 ( .a(n2763), .b(n2764), .out(n1711) );
  xor2 U2341 ( .a(n898), .b(n2765), .out(n2595) );
  xor2 U2342 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[4][0] ), .b(n892), .out(
        n2596) );
  xor2 U2343 ( .a(n2285), .b(\mat_kron/mult_40_G2_G1_G2_G2/ab[2][0] ), .out(
        n2597) );
  xor2 U2344 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[0][7] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[1][6] ), .out(n2766) );
  xor2 U2345 ( .a(n182), .b(\mat_kron/mult_40_G2_G1_G2_G1/ab[2][5] ), .out(
        n2767) );
  xor2 U2346 ( .a(n2766), .b(n2767), .out(n2599) );
  xor2 U2347 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[3][4] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[4][3] ), .out(n2768) );
  xor2 U2348 ( .a(n900), .b(n906), .out(n2769) );
  xor2 U2349 ( .a(n2768), .b(n2769), .out(n2600) );
  xor2 U2350 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[5][2] ), .b(
        \mat_kron/mult_40_G2_G1_G2_G1/ab[6][1] ), .out(n2770) );
  xor2 U2351 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[7][0] ), .b(n915), .out(
        n2771) );
  xor2 U2352 ( .a(n2770), .b(n2771), .out(n1732) );
  xor2 U2353 ( .a(n942), .b(n2772), .out(n2601) );
  xor2 U2354 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[4][0] ), .b(n936), .out(
        n2602) );
  xor2 U2355 ( .a(n2303), .b(\mat_kron/mult_40_G2_G1_G2_G1/ab[2][0] ), .out(
        n2603) );
  xor2 U2356 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[0][7] ), .b(
        \mat_kron/mult_40_G2_G1_G2/ab[1][6] ), .out(n2773) );
  xor2 U2357 ( .a(n177), .b(\mat_kron/mult_40_G2_G1_G2/ab[2][5] ), .out(n2774)
         );
  xor2 U2358 ( .a(n2773), .b(n2774), .out(n2605) );
  xor2 U2359 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[3][4] ), .b(
        \mat_kron/mult_40_G2_G1_G2/ab[4][3] ), .out(n2775) );
  xor2 U2360 ( .a(n944), .b(n950), .out(n2776) );
  xor2 U2361 ( .a(n2775), .b(n2776), .out(n2606) );
  xor2 U2362 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[5][2] ), .b(
        \mat_kron/mult_40_G2_G1_G2/ab[6][1] ), .out(n2777) );
  xor2 U2363 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[7][0] ), .b(n959), .out(n2778)
         );
  xor2 U2364 ( .a(n2777), .b(n2778), .out(n1753) );
  xor2 U2365 ( .a(n986), .b(n2779), .out(n2607) );
  xor2 U2366 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[4][0] ), .b(n980), .out(n2608)
         );
  xor2 U2367 ( .a(n2321), .b(\mat_kron/mult_40_G2_G1_G2/ab[2][0] ), .out(n2609) );
  xor2 U2368 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[0][7] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[1][6] ), .out(n2780) );
  xor2 U2369 ( .a(n178), .b(\mat_kron/mult_40_G2_G1_G1_G2/ab[2][5] ), .out(
        n2781) );
  xor2 U2370 ( .a(n2780), .b(n2781), .out(n2611) );
  xor2 U2371 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[3][4] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[4][3] ), .out(n2782) );
  xor2 U2372 ( .a(n988), .b(n994), .out(n2783) );
  xor2 U2373 ( .a(n2782), .b(n2783), .out(n2612) );
  xor2 U2374 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[5][2] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G2/ab[6][1] ), .out(n2784) );
  xor2 U2375 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[7][0] ), .b(n1003), .out(
        n2785) );
  xor2 U2376 ( .a(n2784), .b(n2785), .out(n1774) );
  xor2 U2377 ( .a(n1030), .b(n2786), .out(n2613) );
  xor2 U2378 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[4][0] ), .b(n1024), .out(
        n2614) );
  xor2 U2379 ( .a(n2339), .b(\mat_kron/mult_40_G2_G1_G1_G2/ab[2][0] ), .out(
        n2615) );
  xor2 U2380 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[0][7] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[1][6] ), .out(n2787) );
  xor2 U2381 ( .a(n186), .b(\mat_kron/mult_40_G2_G1_G1_G1/ab[2][5] ), .out(
        n2788) );
  xor2 U2382 ( .a(n2787), .b(n2788), .out(n2617) );
  xor2 U2383 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[3][4] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[4][3] ), .out(n2789) );
  xor2 U2384 ( .a(n1032), .b(n1038), .out(n2790) );
  xor2 U2385 ( .a(n2789), .b(n2790), .out(n2618) );
  xor2 U2386 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[5][2] ), .b(
        \mat_kron/mult_40_G2_G1_G1_G1/ab[6][1] ), .out(n2791) );
  xor2 U2387 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[7][0] ), .b(n1047), .out(
        n2792) );
  xor2 U2388 ( .a(n2791), .b(n2792), .out(n1795) );
  xor2 U2389 ( .a(n1074), .b(n2793), .out(n2619) );
  xor2 U2390 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[4][0] ), .b(n1068), .out(
        n2620) );
  xor2 U2391 ( .a(n2357), .b(\mat_kron/mult_40_G2_G1_G1_G1/ab[2][0] ), .out(
        n2621) );
  xor2 U2392 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[0][7] ), .b(
        \mat_kron/mult_40_G2_G1_G1/ab[1][6] ), .out(n2794) );
  xor2 U2393 ( .a(n185), .b(\mat_kron/mult_40_G2_G1_G1/ab[2][5] ), .out(n2795)
         );
  xor2 U2394 ( .a(n2794), .b(n2795), .out(n2623) );
  xor2 U2395 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[3][4] ), .b(
        \mat_kron/mult_40_G2_G1_G1/ab[4][3] ), .out(n2796) );
  xor2 U2396 ( .a(n1076), .b(n1082), .out(n2797) );
  xor2 U2397 ( .a(n2796), .b(n2797), .out(n2624) );
  xor2 U2398 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[5][2] ), .b(
        \mat_kron/mult_40_G2_G1_G1/ab[6][1] ), .out(n2798) );
  xor2 U2399 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[7][0] ), .b(n1091), .out(n2799) );
  xor2 U2400 ( .a(n2798), .b(n2799), .out(n1816) );
  xor2 U2401 ( .a(n1118), .b(n2800), .out(n2625) );
  xor2 U2402 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[4][0] ), .b(n1112), .out(n2626) );
  xor2 U2403 ( .a(n2375), .b(\mat_kron/mult_40_G2_G1_G1/ab[2][0] ), .out(n2627) );
  xor2 U2404 ( .a(\mat_kron/mult_40_G2_G1/ab[0][7] ), .b(
        \mat_kron/mult_40_G2_G1/ab[1][6] ), .out(n2801) );
  xor2 U2405 ( .a(n183), .b(\mat_kron/mult_40_G2_G1/ab[2][5] ), .out(n2802) );
  xor2 U2406 ( .a(n2801), .b(n2802), .out(n2629) );
  xor2 U2407 ( .a(\mat_kron/mult_40_G2_G1/ab[3][4] ), .b(
        \mat_kron/mult_40_G2_G1/ab[4][3] ), .out(n2803) );
  xor2 U2408 ( .a(n1120), .b(n1126), .out(n2804) );
  xor2 U2409 ( .a(n2803), .b(n2804), .out(n2630) );
  xor2 U2410 ( .a(\mat_kron/mult_40_G2_G1/ab[5][2] ), .b(
        \mat_kron/mult_40_G2_G1/ab[6][1] ), .out(n2805) );
  xor2 U2411 ( .a(\mat_kron/mult_40_G2_G1/ab[7][0] ), .b(n1135), .out(n2806)
         );
  xor2 U2412 ( .a(n2805), .b(n2806), .out(n1837) );
  xor2 U2413 ( .a(n1162), .b(n2807), .out(n2631) );
  xor2 U2414 ( .a(\mat_kron/mult_40_G2_G1/ab[4][0] ), .b(n1156), .out(n2632)
         );
  xor2 U2415 ( .a(n2393), .b(\mat_kron/mult_40_G2_G1/ab[2][0] ), .out(n2633)
         );
  xor2 U2416 ( .a(\mat_kron/mult_40_G2/ab[0][7] ), .b(
        \mat_kron/mult_40_G2/ab[1][6] ), .out(n2808) );
  xor2 U2417 ( .a(n179), .b(\mat_kron/mult_40_G2/ab[2][5] ), .out(n2809) );
  xor2 U2418 ( .a(n2808), .b(n2809), .out(n2635) );
  xor2 U2419 ( .a(\mat_kron/mult_40_G2/ab[3][4] ), .b(
        \mat_kron/mult_40_G2/ab[4][3] ), .out(n2810) );
  xor2 U2420 ( .a(n1164), .b(n1170), .out(n2811) );
  xor2 U2421 ( .a(n2810), .b(n2811), .out(n2636) );
  xor2 U2422 ( .a(\mat_kron/mult_40_G2/ab[5][2] ), .b(
        \mat_kron/mult_40_G2/ab[6][1] ), .out(n2812) );
  xor2 U2423 ( .a(\mat_kron/mult_40_G2/ab[7][0] ), .b(n1179), .out(n2813) );
  xor2 U2424 ( .a(n2812), .b(n2813), .out(n1858) );
  xor2 U2425 ( .a(n1206), .b(n2814), .out(n2637) );
  xor2 U2426 ( .a(\mat_kron/mult_40_G2/ab[4][0] ), .b(n1200), .out(n2638) );
  xor2 U2427 ( .a(n2411), .b(\mat_kron/mult_40_G2/ab[2][0] ), .out(n2639) );
  xor2 U2428 ( .a(\mat_kron/mult_40/ab[0][7] ), .b(\mat_kron/mult_40/ab[1][6] ), .out(n2815) );
  xor2 U2429 ( .a(n187), .b(\mat_kron/mult_40/ab[2][5] ), .out(n2816) );
  xor2 U2430 ( .a(n2815), .b(n2816), .out(n2641) );
  xor2 U2431 ( .a(\mat_kron/mult_40/ab[3][4] ), .b(\mat_kron/mult_40/ab[4][3] ), .out(n2817) );
  xor2 U2432 ( .a(n1208), .b(n1214), .out(n2818) );
  xor2 U2433 ( .a(n2817), .b(n2818), .out(n2642) );
  xor2 U2434 ( .a(\mat_kron/mult_40/ab[5][2] ), .b(\mat_kron/mult_40/ab[6][1] ), .out(n2819) );
  xor2 U2435 ( .a(\mat_kron/mult_40/ab[7][0] ), .b(n1223), .out(n2820) );
  xor2 U2436 ( .a(n2819), .b(n2820), .out(n1879) );
  xor2 U2437 ( .a(n1250), .b(n2821), .out(n2643) );
  xor2 U2438 ( .a(\mat_kron/mult_40/ab[4][0] ), .b(n1244), .out(n2644) );
  xor2 U2439 ( .a(n2429), .b(\mat_kron/mult_40/ab[2][0] ), .out(n2645) );
  xor2 U2440 ( .a(A[9]), .b(\mat_sub/r102/B_AS [1]), .out(n1882) );
  xor2 U2441 ( .a(A[25]), .b(\mat_sub/r94/B_AS [1]), .out(n1895) );
  xor2 U2442 ( .a(A[1]), .b(\mat_sub/r106/B_AS [1]), .out(n1900) );
  xor2 U2443 ( .a(A[17]), .b(\mat_sub/r98/B_AS [1]), .out(n1903) );
  xor2 U2444 ( .a(n2466), .b(n2822), .out(n2646) );
  xor2 U2445 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[7] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[7] ), .out(n1912) );
  xor2 U2446 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ), .out(n1914) );
  xor2 U2447 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ), .out(n1918) );
  xor2 U2448 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[7] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[7] ), .out(n1923) );
  xor2 U2449 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ), .out(n1925) );
  xor2 U2450 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ), .out(n1927) );
  xor2 U2451 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ), .out(n1931) );
  xor2 U2452 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ), .out(n1935) );
  xor2 U2453 ( .a(n2472), .b(n2823), .out(n2647) );
  xor2 U2454 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[7] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[7] ), .out(n1938) );
  xor2 U2455 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ), .out(n1940) );
  xor2 U2456 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ), .out(n1944) );
  xor2 U2457 ( .a(n2467), .b(n2824), .out(n2648) );
  xor2 U2458 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ), .out(n1948) );
  xor2 U2459 ( .a(n2477), .b(n2825), .out(n2649) );
  xor2 U2460 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[7] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[7] ), .out(n1951) );
  xor2 U2461 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ), .out(n1953) );
  xor2 U2462 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ), .out(n1957) );
  xor2 U2463 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ), .out(n1961) );
  xor2 U2464 ( .a(A[6]), .b(\mat_add/r106/B_AS [6]), .out(n1963) );
  xor2 U2465 ( .a(A[4]), .b(\mat_add/r106/B_AS [4]), .out(n1967) );
  xor2 U2466 ( .a(A[30]), .b(\mat_add/r94/B_AS [6]), .out(n1971) );
  xor2 U2467 ( .a(A[2]), .b(\mat_add/r106/B_AS [2]), .out(n1973) );
  xor2 U2468 ( .a(A[28]), .b(\mat_add/r94/B_AS [4]), .out(n1977) );
  xor2 U2469 ( .a(A[26]), .b(\mat_add/r94/B_AS [2]), .out(n1981) );
  xor2 U2470 ( .a(A[22]), .b(\mat_add/r98/B_AS [6]), .out(n1983) );
  xor2 U2471 ( .a(A[20]), .b(\mat_add/r98/B_AS [4]), .out(n1987) );
  xor2 U2472 ( .a(A[18]), .b(\mat_add/r98/B_AS [2]), .out(n1991) );
  xor2 U2473 ( .a(A[14]), .b(\mat_add/r102/B_AS [6]), .out(n1993) );
  xor2 U2474 ( .a(A[12]), .b(\mat_add/r102/B_AS [4]), .out(n1997) );
  xor2 U2475 ( .a(A[10]), .b(\mat_add/r102/B_AS [2]), .out(n2001) );
  nor2 U2476 ( .a(n199), .b(\mat_mul/mult_37_G2_G2_G2/ab[2][4] ), .out(n2826)
         );
  nor2 U2477 ( .a(n205), .b(\mat_mul/mult_37_G2_G2_G2/ab[3][3] ), .out(n2827)
         );
  inv U2478 ( .in(n2006), .out(n214) );
  nor2 U2479 ( .a(n214), .b(\mat_mul/mult_37_G2_G2_G2/ab[4][2] ), .out(n2828)
         );
  inv U2480 ( .in(n223), .out(n2829) );
  oai22 U2481 ( .a(n2829), .b(n2014), .c(n222), .d(n1387), .out(n2830) );
  nor2 U2482 ( .a(n2660), .b(\mat_mul/mult_37_G2_G2_G2/ab[6][0] ), .out(n237)
         );
  nor2 U2483 ( .a(n287), .b(\mat_mul/mult_37_G2_G2/ab[2][4] ), .out(n2831) );
  nor2 U2484 ( .a(n293), .b(\mat_mul/mult_37_G2_G2/ab[3][3] ), .out(n2832) );
  inv U2485 ( .in(n2042), .out(n302) );
  nor2 U2486 ( .a(n302), .b(\mat_mul/mult_37_G2_G2/ab[4][2] ), .out(n2833) );
  inv U2487 ( .in(n311), .out(n2834) );
  oai22 U2488 ( .a(n2834), .b(n2050), .c(n310), .d(n1429), .out(n2835) );
  nor2 U2489 ( .a(n2674), .b(\mat_mul/mult_37_G2_G2/ab[6][0] ), .out(n325) );
  oai22 U2490 ( .a(n2836), .b(n2824), .c(n1314), .d(n2467), .out(n1926) );
  aoi22 U2491 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ), .c(n1926), .d(n2837), .out(n1920) );
  oai22 U2492 ( .a(n2468), .b(n2469), .c(n1920), .d(n1318), .out(n1917) );
  aoi22 U2493 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ), .c(n1917), .d(n2838), .out(n1916) );
  oai22 U2494 ( .a(n2470), .b(n2471), .c(n1916), .d(n1320), .out(n1913) );
  aoi22 U2495 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ), .c(n1913), .d(n2839), .out(n1911) );
  xor2 U2496 ( .a(n2840), .b(n203), .out(n212) );
  xor2 U2497 ( .a(n2841), .b(n1385), .out(n2018) );
  xor2 U2498 ( .a(n2842), .b(n1382), .out(n1394) );
  xor2 U2499 ( .a(n2843), .b(n1387), .out(n236) );
  xor2 U2500 ( .a(n2844), .b(n291), .out(n300) );
  xor2 U2501 ( .a(n2845), .b(n1427), .out(n2054) );
  xor2 U2502 ( .a(n2846), .b(n1424), .out(n1436) );
  xor2 U2503 ( .a(n2847), .b(n1429), .out(n324) );
  xor2 U2504 ( .a(n201), .b(n2005), .out(n1383) );
  xor2 U2505 ( .a(n199), .b(\mat_mul/mult_37_G2_G2_G2/ab[2][4] ), .out(n1378)
         );
  xor2 U2506 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[3][3] ), .b(n205), .out(n2840)
         );
  xor2 U2507 ( .a(n2002), .b(\mat_mul/mult_37_G2_G2_G2/ab[2][2] ), .out(n1386)
         );
  xor2 U2508 ( .a(n209), .b(n2007), .out(n2842) );
  xor2 U2509 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[4][2] ), .b(n2006), .out(n1388)
         );
  xor2 U2510 ( .a(n217), .b(n216), .out(n1391) );
  xor2 U2511 ( .a(n2011), .b(n219), .out(n2848) );
  xor2 U2512 ( .a(n2012), .b(n221), .out(n1393) );
  xor2 U2513 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[5][1] ), .b(n223), .out(n2843)
         );
  xor2 U2514 ( .a(n2830), .b(n235), .out(n2849) );
  xor2 U2515 ( .a(n2849), .b(n2502), .out(n1395) );
  xor2 U2516 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[5][0] ), .b(n234), .out(n1397)
         );
  xor2 U2517 ( .a(\mat_mul/mult_37_G2_G2_G2/ab[3][0] ), .b(n2016), .out(n1398)
         );
  xor2 U2518 ( .a(n289), .b(n2041), .out(n1425) );
  xor2 U2519 ( .a(n287), .b(\mat_mul/mult_37_G2_G2/ab[2][4] ), .out(n1420) );
  xor2 U2520 ( .a(\mat_mul/mult_37_G2_G2/ab[3][3] ), .b(n293), .out(n2844) );
  xor2 U2521 ( .a(n2038), .b(\mat_mul/mult_37_G2_G2/ab[2][2] ), .out(n1428) );
  xor2 U2522 ( .a(n297), .b(n2043), .out(n2846) );
  xor2 U2523 ( .a(\mat_mul/mult_37_G2_G2/ab[4][2] ), .b(n2042), .out(n1430) );
  xor2 U2524 ( .a(n305), .b(n304), .out(n1433) );
  xor2 U2525 ( .a(n2047), .b(n307), .out(n2850) );
  xor2 U2526 ( .a(n2048), .b(n309), .out(n1435) );
  xor2 U2527 ( .a(\mat_mul/mult_37_G2_G2/ab[5][1] ), .b(n311), .out(n2847) );
  xor2 U2528 ( .a(n2835), .b(n323), .out(n2851) );
  xor2 U2529 ( .a(n2851), .b(n2514), .out(n1437) );
  xor2 U2530 ( .a(\mat_mul/mult_37_G2_G2/ab[5][0] ), .b(n322), .out(n1439) );
  xor2 U2531 ( .a(\mat_mul/mult_37_G2_G2/ab[3][0] ), .b(n2052), .out(n1440) );
  xor2 U2532 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ), .b(n2471), .out(n1915) );
  xor2 U2533 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ), .b(n2469), .out(n1919) );
  nor2 U2534 ( .a(n243), .b(\mat_mul/mult_37_G2_G2_G1/ab[2][4] ), .out(n2852)
         );
  nor2 U2535 ( .a(n249), .b(\mat_mul/mult_37_G2_G2_G1/ab[3][3] ), .out(n2853)
         );
  inv U2536 ( .in(n2024), .out(n258) );
  nor2 U2537 ( .a(n258), .b(\mat_mul/mult_37_G2_G2_G1/ab[4][2] ), .out(n2854)
         );
  inv U2538 ( .in(n267), .out(n2855) );
  oai22 U2539 ( .a(n2855), .b(n2032), .c(n266), .d(n1408), .out(n2856) );
  nor2 U2540 ( .a(n2667), .b(\mat_mul/mult_37_G2_G2_G1/ab[6][0] ), .out(n281)
         );
  nor2 U2541 ( .a(n419), .b(\mat_mul/mult_37_G2_G1/ab[2][4] ), .out(n2857) );
  nor2 U2542 ( .a(n425), .b(\mat_mul/mult_37_G2_G1/ab[3][3] ), .out(n2858) );
  inv U2543 ( .in(n2096), .out(n434) );
  nor2 U2544 ( .a(n434), .b(\mat_mul/mult_37_G2_G1/ab[4][2] ), .out(n2859) );
  inv U2545 ( .in(n443), .out(n2860) );
  oai22 U2546 ( .a(n2860), .b(n2104), .c(n442), .d(n1492), .out(n2861) );
  nor2 U2547 ( .a(n2695), .b(\mat_mul/mult_37_G2_G1/ab[6][0] ), .out(n457) );
  oai22 U2548 ( .a(n2862), .b(n2825), .c(n1330), .d(n2477), .out(n1947) );
  aoi22 U2549 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ), .c(n1947), .d(n2863), .out(n1946) );
  oai22 U2550 ( .a(n2478), .b(n2479), .c(n1946), .d(n1334), .out(n1943) );
  aoi22 U2551 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ), .c(n1943), .d(n2864), .out(n1942) );
  oai22 U2552 ( .a(n2480), .b(n2481), .c(n1942), .d(n1336), .out(n1939) );
  aoi22 U2553 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ), .c(n1939), .d(n2865), .out(n1937) );
  xor2 U2554 ( .a(n2866), .b(n247), .out(n256) );
  xor2 U2555 ( .a(n2867), .b(n1406), .out(n2036) );
  xor2 U2556 ( .a(n2868), .b(n1403), .out(n1415) );
  xor2 U2557 ( .a(n2869), .b(n1408), .out(n280) );
  xor2 U2558 ( .a(n2870), .b(n423), .out(n432) );
  xor2 U2559 ( .a(n2871), .b(n1490), .out(n2108) );
  xor2 U2560 ( .a(n2872), .b(n1487), .out(n1499) );
  xor2 U2561 ( .a(n2873), .b(n1492), .out(n456) );
  xor2 U2562 ( .a(n245), .b(n2023), .out(n1404) );
  xor2 U2563 ( .a(n243), .b(\mat_mul/mult_37_G2_G2_G1/ab[2][4] ), .out(n1399)
         );
  xor2 U2564 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[3][3] ), .b(n249), .out(n2866)
         );
  xor2 U2565 ( .a(n2020), .b(\mat_mul/mult_37_G2_G2_G1/ab[2][2] ), .out(n1407)
         );
  xor2 U2566 ( .a(n253), .b(n2025), .out(n2868) );
  xor2 U2567 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[4][2] ), .b(n2024), .out(n1409)
         );
  xor2 U2568 ( .a(n261), .b(n260), .out(n1412) );
  xor2 U2569 ( .a(n2029), .b(n263), .out(n2874) );
  xor2 U2570 ( .a(n2030), .b(n265), .out(n1414) );
  xor2 U2571 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[5][1] ), .b(n267), .out(n2869)
         );
  xor2 U2572 ( .a(n2856), .b(n279), .out(n2875) );
  xor2 U2573 ( .a(n2875), .b(n2508), .out(n1416) );
  xor2 U2574 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[5][0] ), .b(n278), .out(n1418)
         );
  xor2 U2575 ( .a(\mat_mul/mult_37_G2_G2_G1/ab[3][0] ), .b(n2034), .out(n1419)
         );
  xor2 U2576 ( .a(n421), .b(n2095), .out(n1488) );
  xor2 U2577 ( .a(n419), .b(\mat_mul/mult_37_G2_G1/ab[2][4] ), .out(n1483) );
  xor2 U2578 ( .a(\mat_mul/mult_37_G2_G1/ab[3][3] ), .b(n425), .out(n2870) );
  xor2 U2579 ( .a(n2092), .b(\mat_mul/mult_37_G2_G1/ab[2][2] ), .out(n1491) );
  xor2 U2580 ( .a(n429), .b(n2097), .out(n2872) );
  xor2 U2581 ( .a(\mat_mul/mult_37_G2_G1/ab[4][2] ), .b(n2096), .out(n1493) );
  xor2 U2582 ( .a(n437), .b(n436), .out(n1496) );
  xor2 U2583 ( .a(n2101), .b(n439), .out(n2876) );
  xor2 U2584 ( .a(n2102), .b(n441), .out(n1498) );
  xor2 U2585 ( .a(\mat_mul/mult_37_G2_G1/ab[5][1] ), .b(n443), .out(n2873) );
  xor2 U2586 ( .a(n2861), .b(n455), .out(n2877) );
  xor2 U2587 ( .a(n2877), .b(n2532), .out(n1500) );
  xor2 U2588 ( .a(\mat_mul/mult_37_G2_G1/ab[5][0] ), .b(n454), .out(n1502) );
  xor2 U2589 ( .a(\mat_mul/mult_37_G2_G1/ab[3][0] ), .b(n2106), .out(n1503) );
  xor2 U2590 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ), .b(n2481), .out(n1941) );
  xor2 U2591 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ), .b(n2479), .out(n1945) );
  nor2 U2592 ( .a(n331), .b(\mat_mul/mult_37_G2_G1_G2/ab[2][4] ), .out(n2878)
         );
  nor2 U2593 ( .a(n337), .b(\mat_mul/mult_37_G2_G1_G2/ab[3][3] ), .out(n2879)
         );
  inv U2594 ( .in(n2060), .out(n346) );
  nor2 U2595 ( .a(n346), .b(\mat_mul/mult_37_G2_G1_G2/ab[4][2] ), .out(n2880)
         );
  inv U2596 ( .in(n355), .out(n2881) );
  oai22 U2597 ( .a(n2881), .b(n2068), .c(n354), .d(n1450), .out(n2882) );
  nor2 U2598 ( .a(n2681), .b(\mat_mul/mult_37_G2_G1_G2/ab[6][0] ), .out(n369)
         );
  nor2 U2599 ( .a(n463), .b(\mat_mul/mult_37_G2/ab[2][4] ), .out(n2883) );
  nor2 U2600 ( .a(n469), .b(\mat_mul/mult_37_G2/ab[3][3] ), .out(n2884) );
  inv U2601 ( .in(n2114), .out(n478) );
  nor2 U2602 ( .a(n478), .b(\mat_mul/mult_37_G2/ab[4][2] ), .out(n2885) );
  inv U2603 ( .in(n487), .out(n2886) );
  oai22 U2604 ( .a(n2886), .b(n2122), .c(n486), .d(n1513), .out(n2887) );
  nor2 U2605 ( .a(n2702), .b(\mat_mul/mult_37_G2/ab[6][0] ), .out(n501) );
  oai22 U2606 ( .a(n2822), .b(n2888), .c(n1338), .d(n2466), .out(n1960) );
  aoi22 U2607 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ), .c(n1960), .d(n2889), .out(n1959) );
  oai22 U2608 ( .a(n2482), .b(n2483), .c(n1959), .d(n1342), .out(n1956) );
  aoi22 U2609 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ), .c(n1956), .d(n2890), .out(n1955) );
  oai22 U2610 ( .a(n2484), .b(n2485), .c(n1955), .d(n1344), .out(n1952) );
  aoi22 U2611 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ), .c(n1952), .d(n2891), .out(n1950) );
  xor2 U2612 ( .a(n2892), .b(n335), .out(n344) );
  xor2 U2613 ( .a(n2893), .b(n1448), .out(n2072) );
  xor2 U2614 ( .a(n2894), .b(n1445), .out(n1457) );
  xor2 U2615 ( .a(n2895), .b(n1450), .out(n368) );
  xor2 U2616 ( .a(n2896), .b(n467), .out(n476) );
  xor2 U2617 ( .a(n2897), .b(n1511), .out(n2126) );
  xor2 U2618 ( .a(n2898), .b(n1508), .out(n1520) );
  xor2 U2619 ( .a(n2899), .b(n1513), .out(n500) );
  inv U2620 ( .in(n1340), .out(n2822) );
  inv U2621 ( .in(n1339), .out(n2888) );
  xor2 U2622 ( .a(n333), .b(n2059), .out(n1446) );
  xor2 U2623 ( .a(n331), .b(\mat_mul/mult_37_G2_G1_G2/ab[2][4] ), .out(n1441)
         );
  xor2 U2624 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[3][3] ), .b(n337), .out(n2892)
         );
  xor2 U2625 ( .a(n2056), .b(\mat_mul/mult_37_G2_G1_G2/ab[2][2] ), .out(n1449)
         );
  xor2 U2626 ( .a(n341), .b(n2061), .out(n2894) );
  xor2 U2627 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[4][2] ), .b(n2060), .out(n1451)
         );
  xor2 U2628 ( .a(n349), .b(n348), .out(n1454) );
  xor2 U2629 ( .a(n2065), .b(n351), .out(n2900) );
  xor2 U2630 ( .a(n2066), .b(n353), .out(n1456) );
  xor2 U2631 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[5][1] ), .b(n355), .out(n2895)
         );
  xor2 U2632 ( .a(n2882), .b(n367), .out(n2901) );
  xor2 U2633 ( .a(n2901), .b(n2520), .out(n1458) );
  xor2 U2634 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[5][0] ), .b(n366), .out(n1460)
         );
  xor2 U2635 ( .a(\mat_mul/mult_37_G2_G1_G2/ab[3][0] ), .b(n2070), .out(n1461)
         );
  xor2 U2636 ( .a(n465), .b(n2113), .out(n1509) );
  xor2 U2637 ( .a(n463), .b(\mat_mul/mult_37_G2/ab[2][4] ), .out(n1504) );
  xor2 U2638 ( .a(\mat_mul/mult_37_G2/ab[3][3] ), .b(n469), .out(n2896) );
  xor2 U2639 ( .a(n2110), .b(\mat_mul/mult_37_G2/ab[2][2] ), .out(n1512) );
  xor2 U2640 ( .a(n473), .b(n2115), .out(n2898) );
  xor2 U2641 ( .a(\mat_mul/mult_37_G2/ab[4][2] ), .b(n2114), .out(n1514) );
  xor2 U2642 ( .a(n481), .b(n480), .out(n1517) );
  xor2 U2643 ( .a(n2119), .b(n483), .out(n2902) );
  xor2 U2644 ( .a(n2120), .b(n485), .out(n1519) );
  xor2 U2645 ( .a(\mat_mul/mult_37_G2/ab[5][1] ), .b(n487), .out(n2899) );
  xor2 U2646 ( .a(n2887), .b(n499), .out(n2903) );
  xor2 U2647 ( .a(n2903), .b(n2538), .out(n1521) );
  xor2 U2648 ( .a(\mat_mul/mult_37_G2/ab[5][0] ), .b(n498), .out(n1523) );
  xor2 U2649 ( .a(\mat_mul/mult_37_G2/ab[3][0] ), .b(n2124), .out(n1524) );
  xor2 U2650 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ), .b(n2485), .out(n1954) );
  xor2 U2651 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ), .b(n2483), .out(n1958) );
  nor2 U2652 ( .a(n375), .b(\mat_mul/mult_37_G2_G1_G1/ab[2][4] ), .out(n2904)
         );
  nor2 U2653 ( .a(n381), .b(\mat_mul/mult_37_G2_G1_G1/ab[3][3] ), .out(n2905)
         );
  inv U2654 ( .in(n2078), .out(n390) );
  nor2 U2655 ( .a(n390), .b(\mat_mul/mult_37_G2_G1_G1/ab[4][2] ), .out(n2906)
         );
  inv U2656 ( .in(n399), .out(n2907) );
  oai22 U2657 ( .a(n2907), .b(n2086), .c(n398), .d(n1471), .out(n2908) );
  nor2 U2658 ( .a(n2688), .b(\mat_mul/mult_37_G2_G1_G1/ab[6][0] ), .out(n413)
         );
  nor2 U2659 ( .a(n507), .b(\mat_mul/mult_37/ab[2][4] ), .out(n2909) );
  nor2 U2660 ( .a(n513), .b(\mat_mul/mult_37/ab[3][3] ), .out(n2910) );
  inv U2661 ( .in(n2132), .out(n522) );
  nor2 U2662 ( .a(n522), .b(\mat_mul/mult_37/ab[4][2] ), .out(n2911) );
  inv U2663 ( .in(n531), .out(n2912) );
  oai22 U2664 ( .a(n2912), .b(n2140), .c(n530), .d(n1534), .out(n2913) );
  nor2 U2665 ( .a(n2709), .b(\mat_mul/mult_37/ab[6][0] ), .out(n545) );
  oai22 U2666 ( .a(n2914), .b(n2823), .c(n1322), .d(n2472), .out(n1934) );
  aoi22 U2667 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ), .c(n1934), .d(n2915), .out(n1933) );
  oai22 U2668 ( .a(n2473), .b(n2474), .c(n1933), .d(n1326), .out(n1930) );
  aoi22 U2669 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ), .c(n1930), .d(n2916), .out(n1929) );
  oai22 U2670 ( .a(n2475), .b(n2476), .c(n1929), .d(n1328), .out(n1924) );
  aoi22 U2671 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ), .b(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ), .c(n1924), .d(n2917), .out(n1922) );
  xor2 U2672 ( .a(n2918), .b(n379), .out(n388) );
  xor2 U2673 ( .a(n2919), .b(n1469), .out(n2090) );
  xor2 U2674 ( .a(n2920), .b(n1466), .out(n1478) );
  xor2 U2675 ( .a(n2921), .b(n1471), .out(n412) );
  xor2 U2676 ( .a(n2922), .b(n511), .out(n520) );
  xor2 U2677 ( .a(n2923), .b(n1532), .out(n2144) );
  xor2 U2678 ( .a(n2924), .b(n1529), .out(n1541) );
  xor2 U2679 ( .a(n2925), .b(n1534), .out(n544) );
  xor2 U2680 ( .a(n377), .b(n2077), .out(n1467) );
  xor2 U2681 ( .a(n375), .b(\mat_mul/mult_37_G2_G1_G1/ab[2][4] ), .out(n1462)
         );
  xor2 U2682 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[3][3] ), .b(n381), .out(n2918)
         );
  xor2 U2683 ( .a(n2074), .b(\mat_mul/mult_37_G2_G1_G1/ab[2][2] ), .out(n1470)
         );
  xor2 U2684 ( .a(n385), .b(n2079), .out(n2920) );
  xor2 U2685 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[4][2] ), .b(n2078), .out(n1472)
         );
  xor2 U2686 ( .a(n393), .b(n392), .out(n1475) );
  xor2 U2687 ( .a(n2083), .b(n395), .out(n2926) );
  xor2 U2688 ( .a(n2084), .b(n397), .out(n1477) );
  xor2 U2689 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[5][1] ), .b(n399), .out(n2921)
         );
  xor2 U2690 ( .a(n2908), .b(n411), .out(n2927) );
  xor2 U2691 ( .a(n2927), .b(n2526), .out(n1479) );
  xor2 U2692 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[5][0] ), .b(n410), .out(n1481)
         );
  xor2 U2693 ( .a(\mat_mul/mult_37_G2_G1_G1/ab[3][0] ), .b(n2088), .out(n1482)
         );
  xor2 U2694 ( .a(n509), .b(n2131), .out(n1530) );
  xor2 U2695 ( .a(n507), .b(\mat_mul/mult_37/ab[2][4] ), .out(n1525) );
  xor2 U2696 ( .a(\mat_mul/mult_37/ab[3][3] ), .b(n513), .out(n2922) );
  xor2 U2697 ( .a(n2128), .b(\mat_mul/mult_37/ab[2][2] ), .out(n1533) );
  xor2 U2698 ( .a(n517), .b(n2133), .out(n2924) );
  xor2 U2699 ( .a(\mat_mul/mult_37/ab[4][2] ), .b(n2132), .out(n1535) );
  xor2 U2700 ( .a(n525), .b(n524), .out(n1538) );
  xor2 U2701 ( .a(n2137), .b(n527), .out(n2928) );
  xor2 U2702 ( .a(n2138), .b(n529), .out(n1540) );
  xor2 U2703 ( .a(\mat_mul/mult_37/ab[5][1] ), .b(n531), .out(n2925) );
  xor2 U2704 ( .a(n2913), .b(n543), .out(n2929) );
  xor2 U2705 ( .a(n2929), .b(n2544), .out(n1542) );
  xor2 U2706 ( .a(\mat_mul/mult_37/ab[5][0] ), .b(n542), .out(n1544) );
  xor2 U2707 ( .a(\mat_mul/mult_37/ab[3][0] ), .b(n2142), .out(n1545) );
  xor2 U2708 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ), .b(n2476), .out(n1928) );
  xor2 U2709 ( .a(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ), .b(n2474), .out(n1932) );
  nor2 U2710 ( .a(n551), .b(\mat_kron/mult_40_G2_G2_G2_G2/ab[2][4] ), .out(
        n2930) );
  nor2 U2711 ( .a(n557), .b(\mat_kron/mult_40_G2_G2_G2_G2/ab[3][3] ), .out(
        n2931) );
  inv U2712 ( .in(n2150), .out(n566) );
  nor2 U2713 ( .a(n566), .b(\mat_kron/mult_40_G2_G2_G2_G2/ab[4][2] ), .out(
        n2932) );
  inv U2714 ( .in(n575), .out(n2933) );
  oai22 U2715 ( .a(n2933), .b(n2158), .c(n574), .d(n1555), .out(n2934) );
  nor2 U2716 ( .a(n2716), .b(\mat_kron/mult_40_G2_G2_G2_G2/ab[6][0] ), .out(
        n589) );
  xor2 U2717 ( .a(n2935), .b(n555), .out(n564) );
  xor2 U2718 ( .a(n2936), .b(n1553), .out(n2162) );
  xor2 U2719 ( .a(n2937), .b(n1550), .out(n1562) );
  xor2 U2720 ( .a(n2938), .b(n1555), .out(n588) );
  xor2 U2721 ( .a(n553), .b(n2149), .out(n1551) );
  xor2 U2722 ( .a(n551), .b(\mat_kron/mult_40_G2_G2_G2_G2/ab[2][4] ), .out(
        n1546) );
  xor2 U2723 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[3][3] ), .b(n557), .out(
        n2935) );
  xor2 U2724 ( .a(n2146), .b(\mat_kron/mult_40_G2_G2_G2_G2/ab[2][2] ), .out(
        n1554) );
  xor2 U2725 ( .a(n561), .b(n2151), .out(n2937) );
  xor2 U2726 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[4][2] ), .b(n2150), .out(
        n1556) );
  xor2 U2727 ( .a(n569), .b(n568), .out(n1559) );
  xor2 U2728 ( .a(n2155), .b(n571), .out(n2939) );
  xor2 U2729 ( .a(n2156), .b(n573), .out(n1561) );
  xor2 U2730 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[5][1] ), .b(n575), .out(
        n2938) );
  xor2 U2731 ( .a(n2934), .b(n587), .out(n2940) );
  xor2 U2732 ( .a(n2940), .b(n2550), .out(n1563) );
  xor2 U2733 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[5][0] ), .b(n586), .out(
        n1565) );
  xor2 U2734 ( .a(\mat_kron/mult_40_G2_G2_G2_G2/ab[3][0] ), .b(n2160), .out(
        n1566) );
  nor2 U2735 ( .a(n595), .b(\mat_kron/mult_40_G2_G2_G2_G1/ab[2][4] ), .out(
        n2941) );
  nor2 U2736 ( .a(n601), .b(\mat_kron/mult_40_G2_G2_G2_G1/ab[3][3] ), .out(
        n2942) );
  inv U2737 ( .in(n2168), .out(n610) );
  nor2 U2738 ( .a(n610), .b(\mat_kron/mult_40_G2_G2_G2_G1/ab[4][2] ), .out(
        n2943) );
  inv U2739 ( .in(n619), .out(n2944) );
  oai22 U2740 ( .a(n2944), .b(n2176), .c(n618), .d(n1576), .out(n2945) );
  nor2 U2741 ( .a(n2723), .b(\mat_kron/mult_40_G2_G2_G2_G1/ab[6][0] ), .out(
        n633) );
  xor2 U2742 ( .a(n2946), .b(n599), .out(n608) );
  xor2 U2743 ( .a(n2947), .b(n1574), .out(n2180) );
  xor2 U2744 ( .a(n2948), .b(n1571), .out(n1583) );
  xor2 U2745 ( .a(n2949), .b(n1576), .out(n632) );
  xor2 U2746 ( .a(n597), .b(n2167), .out(n1572) );
  xor2 U2747 ( .a(n595), .b(\mat_kron/mult_40_G2_G2_G2_G1/ab[2][4] ), .out(
        n1567) );
  xor2 U2748 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[3][3] ), .b(n601), .out(
        n2946) );
  xor2 U2749 ( .a(n2164), .b(\mat_kron/mult_40_G2_G2_G2_G1/ab[2][2] ), .out(
        n1575) );
  xor2 U2750 ( .a(n605), .b(n2169), .out(n2948) );
  xor2 U2751 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[4][2] ), .b(n2168), .out(
        n1577) );
  xor2 U2752 ( .a(n613), .b(n612), .out(n1580) );
  xor2 U2753 ( .a(n2173), .b(n615), .out(n2950) );
  xor2 U2754 ( .a(n2174), .b(n617), .out(n1582) );
  xor2 U2755 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[5][1] ), .b(n619), .out(
        n2949) );
  xor2 U2756 ( .a(n2945), .b(n631), .out(n2951) );
  xor2 U2757 ( .a(n2951), .b(n2556), .out(n1584) );
  xor2 U2758 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[5][0] ), .b(n630), .out(
        n1586) );
  xor2 U2759 ( .a(\mat_kron/mult_40_G2_G2_G2_G1/ab[3][0] ), .b(n2178), .out(
        n1587) );
  nor2 U2760 ( .a(n639), .b(\mat_kron/mult_40_G2_G2_G2/ab[2][4] ), .out(n2952)
         );
  nor2 U2761 ( .a(n645), .b(\mat_kron/mult_40_G2_G2_G2/ab[3][3] ), .out(n2953)
         );
  inv U2762 ( .in(n2186), .out(n654) );
  nor2 U2763 ( .a(n654), .b(\mat_kron/mult_40_G2_G2_G2/ab[4][2] ), .out(n2954)
         );
  inv U2764 ( .in(n663), .out(n2955) );
  oai22 U2765 ( .a(n2955), .b(n2194), .c(n662), .d(n1597), .out(n2956) );
  nor2 U2766 ( .a(n2730), .b(\mat_kron/mult_40_G2_G2_G2/ab[6][0] ), .out(n677)
         );
  xor2 U2767 ( .a(n2957), .b(n643), .out(n652) );
  xor2 U2768 ( .a(n2958), .b(n1595), .out(n2198) );
  xor2 U2769 ( .a(n2959), .b(n1592), .out(n1604) );
  xor2 U2770 ( .a(n2960), .b(n1597), .out(n676) );
  xor2 U2771 ( .a(n641), .b(n2185), .out(n1593) );
  xor2 U2772 ( .a(n639), .b(\mat_kron/mult_40_G2_G2_G2/ab[2][4] ), .out(n1588)
         );
  xor2 U2773 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[3][3] ), .b(n645), .out(n2957)
         );
  xor2 U2774 ( .a(n2182), .b(\mat_kron/mult_40_G2_G2_G2/ab[2][2] ), .out(n1596) );
  xor2 U2775 ( .a(n649), .b(n2187), .out(n2959) );
  xor2 U2776 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[4][2] ), .b(n2186), .out(n1598) );
  xor2 U2777 ( .a(n657), .b(n656), .out(n1601) );
  xor2 U2778 ( .a(n2191), .b(n659), .out(n2961) );
  xor2 U2779 ( .a(n2192), .b(n661), .out(n1603) );
  xor2 U2780 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[5][1] ), .b(n663), .out(n2960)
         );
  xor2 U2781 ( .a(n2956), .b(n675), .out(n2962) );
  xor2 U2782 ( .a(n2962), .b(n2562), .out(n1605) );
  xor2 U2783 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[5][0] ), .b(n674), .out(n1607)
         );
  xor2 U2784 ( .a(\mat_kron/mult_40_G2_G2_G2/ab[3][0] ), .b(n2196), .out(n1608) );
  nor2 U2785 ( .a(n683), .b(\mat_kron/mult_40_G2_G2_G1_G2/ab[2][4] ), .out(
        n2963) );
  nor2 U2786 ( .a(n689), .b(\mat_kron/mult_40_G2_G2_G1_G2/ab[3][3] ), .out(
        n2964) );
  inv U2787 ( .in(n2204), .out(n698) );
  nor2 U2788 ( .a(n698), .b(\mat_kron/mult_40_G2_G2_G1_G2/ab[4][2] ), .out(
        n2965) );
  inv U2789 ( .in(n707), .out(n2966) );
  oai22 U2790 ( .a(n2966), .b(n2212), .c(n706), .d(n1618), .out(n2967) );
  nor2 U2791 ( .a(n2737), .b(\mat_kron/mult_40_G2_G2_G1_G2/ab[6][0] ), .out(
        n721) );
  xor2 U2792 ( .a(n2968), .b(n687), .out(n696) );
  xor2 U2793 ( .a(n2969), .b(n1616), .out(n2216) );
  xor2 U2794 ( .a(n2970), .b(n1613), .out(n1625) );
  xor2 U2795 ( .a(n2971), .b(n1618), .out(n720) );
  xor2 U2796 ( .a(n685), .b(n2203), .out(n1614) );
  xor2 U2797 ( .a(n683), .b(\mat_kron/mult_40_G2_G2_G1_G2/ab[2][4] ), .out(
        n1609) );
  xor2 U2798 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[3][3] ), .b(n689), .out(
        n2968) );
  xor2 U2799 ( .a(n2200), .b(\mat_kron/mult_40_G2_G2_G1_G2/ab[2][2] ), .out(
        n1617) );
  xor2 U2800 ( .a(n693), .b(n2205), .out(n2970) );
  xor2 U2801 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[4][2] ), .b(n2204), .out(
        n1619) );
  xor2 U2802 ( .a(n701), .b(n700), .out(n1622) );
  xor2 U2803 ( .a(n2209), .b(n703), .out(n2972) );
  xor2 U2804 ( .a(n2210), .b(n705), .out(n1624) );
  xor2 U2805 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[5][1] ), .b(n707), .out(
        n2971) );
  xor2 U2806 ( .a(n2967), .b(n719), .out(n2973) );
  xor2 U2807 ( .a(n2973), .b(n2568), .out(n1626) );
  xor2 U2808 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[5][0] ), .b(n718), .out(
        n1628) );
  xor2 U2809 ( .a(\mat_kron/mult_40_G2_G2_G1_G2/ab[3][0] ), .b(n2214), .out(
        n1629) );
  nor2 U2810 ( .a(n727), .b(\mat_kron/mult_40_G2_G2_G1_G1/ab[2][4] ), .out(
        n2974) );
  nor2 U2811 ( .a(n733), .b(\mat_kron/mult_40_G2_G2_G1_G1/ab[3][3] ), .out(
        n2975) );
  inv U2812 ( .in(n2222), .out(n742) );
  nor2 U2813 ( .a(n742), .b(\mat_kron/mult_40_G2_G2_G1_G1/ab[4][2] ), .out(
        n2976) );
  inv U2814 ( .in(n751), .out(n2977) );
  oai22 U2815 ( .a(n2977), .b(n2230), .c(n750), .d(n1639), .out(n2978) );
  nor2 U2816 ( .a(n2744), .b(\mat_kron/mult_40_G2_G2_G1_G1/ab[6][0] ), .out(
        n765) );
  xor2 U2817 ( .a(n2979), .b(n731), .out(n740) );
  xor2 U2818 ( .a(n2980), .b(n1637), .out(n2234) );
  xor2 U2819 ( .a(n2981), .b(n1634), .out(n1646) );
  xor2 U2820 ( .a(n2982), .b(n1639), .out(n764) );
  xor2 U2821 ( .a(n729), .b(n2221), .out(n1635) );
  xor2 U2822 ( .a(n727), .b(\mat_kron/mult_40_G2_G2_G1_G1/ab[2][4] ), .out(
        n1630) );
  xor2 U2823 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[3][3] ), .b(n733), .out(
        n2979) );
  xor2 U2824 ( .a(n2218), .b(\mat_kron/mult_40_G2_G2_G1_G1/ab[2][2] ), .out(
        n1638) );
  xor2 U2825 ( .a(n737), .b(n2223), .out(n2981) );
  xor2 U2826 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[4][2] ), .b(n2222), .out(
        n1640) );
  xor2 U2827 ( .a(n745), .b(n744), .out(n1643) );
  xor2 U2828 ( .a(n2227), .b(n747), .out(n2983) );
  xor2 U2829 ( .a(n2228), .b(n749), .out(n1645) );
  xor2 U2830 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[5][1] ), .b(n751), .out(
        n2982) );
  xor2 U2831 ( .a(n2978), .b(n763), .out(n2984) );
  xor2 U2832 ( .a(n2984), .b(n2574), .out(n1647) );
  xor2 U2833 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[5][0] ), .b(n762), .out(
        n1649) );
  xor2 U2834 ( .a(\mat_kron/mult_40_G2_G2_G1_G1/ab[3][0] ), .b(n2232), .out(
        n1650) );
  nor2 U2835 ( .a(n771), .b(\mat_kron/mult_40_G2_G2_G1/ab[2][4] ), .out(n2985)
         );
  nor2 U2836 ( .a(n777), .b(\mat_kron/mult_40_G2_G2_G1/ab[3][3] ), .out(n2986)
         );
  inv U2837 ( .in(n2240), .out(n786) );
  nor2 U2838 ( .a(n786), .b(\mat_kron/mult_40_G2_G2_G1/ab[4][2] ), .out(n2987)
         );
  inv U2839 ( .in(n795), .out(n2988) );
  oai22 U2840 ( .a(n2988), .b(n2248), .c(n794), .d(n1660), .out(n2989) );
  nor2 U2841 ( .a(n2751), .b(\mat_kron/mult_40_G2_G2_G1/ab[6][0] ), .out(n809)
         );
  xor2 U2842 ( .a(n2990), .b(n775), .out(n784) );
  xor2 U2843 ( .a(n2991), .b(n1658), .out(n2252) );
  xor2 U2844 ( .a(n2992), .b(n1655), .out(n1667) );
  xor2 U2845 ( .a(n2993), .b(n1660), .out(n808) );
  xor2 U2846 ( .a(n773), .b(n2239), .out(n1656) );
  xor2 U2847 ( .a(n771), .b(\mat_kron/mult_40_G2_G2_G1/ab[2][4] ), .out(n1651)
         );
  xor2 U2848 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[3][3] ), .b(n777), .out(n2990)
         );
  xor2 U2849 ( .a(n2236), .b(\mat_kron/mult_40_G2_G2_G1/ab[2][2] ), .out(n1659) );
  xor2 U2850 ( .a(n781), .b(n2241), .out(n2992) );
  xor2 U2851 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[4][2] ), .b(n2240), .out(n1661) );
  xor2 U2852 ( .a(n789), .b(n788), .out(n1664) );
  xor2 U2853 ( .a(n2245), .b(n791), .out(n2994) );
  xor2 U2854 ( .a(n2246), .b(n793), .out(n1666) );
  xor2 U2855 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[5][1] ), .b(n795), .out(n2993)
         );
  xor2 U2856 ( .a(n2989), .b(n807), .out(n2995) );
  xor2 U2857 ( .a(n2995), .b(n2580), .out(n1668) );
  xor2 U2858 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[5][0] ), .b(n806), .out(n1670)
         );
  xor2 U2859 ( .a(\mat_kron/mult_40_G2_G2_G1/ab[3][0] ), .b(n2250), .out(n1671) );
  nor2 U2860 ( .a(n815), .b(\mat_kron/mult_40_G2_G2/ab[2][4] ), .out(n2996) );
  nor2 U2861 ( .a(n821), .b(\mat_kron/mult_40_G2_G2/ab[3][3] ), .out(n2997) );
  inv U2862 ( .in(n2258), .out(n830) );
  nor2 U2863 ( .a(n830), .b(\mat_kron/mult_40_G2_G2/ab[4][2] ), .out(n2998) );
  inv U2864 ( .in(n839), .out(n2999) );
  oai22 U2865 ( .a(n2999), .b(n2266), .c(n838), .d(n1681), .out(n3000) );
  nor2 U2866 ( .a(n2758), .b(\mat_kron/mult_40_G2_G2/ab[6][0] ), .out(n853) );
  xor2 U2867 ( .a(n3001), .b(n819), .out(n828) );
  xor2 U2868 ( .a(n3002), .b(n1679), .out(n2270) );
  xor2 U2869 ( .a(n3003), .b(n1676), .out(n1688) );
  xor2 U2870 ( .a(n3004), .b(n1681), .out(n852) );
  xor2 U2871 ( .a(n817), .b(n2257), .out(n1677) );
  xor2 U2872 ( .a(n815), .b(\mat_kron/mult_40_G2_G2/ab[2][4] ), .out(n1672) );
  xor2 U2873 ( .a(\mat_kron/mult_40_G2_G2/ab[3][3] ), .b(n821), .out(n3001) );
  xor2 U2874 ( .a(n2254), .b(\mat_kron/mult_40_G2_G2/ab[2][2] ), .out(n1680)
         );
  xor2 U2875 ( .a(n825), .b(n2259), .out(n3003) );
  xor2 U2876 ( .a(\mat_kron/mult_40_G2_G2/ab[4][2] ), .b(n2258), .out(n1682)
         );
  xor2 U2877 ( .a(n833), .b(n832), .out(n1685) );
  xor2 U2878 ( .a(n2263), .b(n835), .out(n3005) );
  xor2 U2879 ( .a(n2264), .b(n837), .out(n1687) );
  xor2 U2880 ( .a(\mat_kron/mult_40_G2_G2/ab[5][1] ), .b(n839), .out(n3004) );
  xor2 U2881 ( .a(n3000), .b(n851), .out(n3006) );
  xor2 U2882 ( .a(n3006), .b(n2586), .out(n1689) );
  xor2 U2883 ( .a(\mat_kron/mult_40_G2_G2/ab[5][0] ), .b(n850), .out(n1691) );
  xor2 U2884 ( .a(\mat_kron/mult_40_G2_G2/ab[3][0] ), .b(n2268), .out(n1692)
         );
  nor2 U2885 ( .a(n859), .b(\mat_kron/mult_40_G2_G1_G2_G2/ab[2][4] ), .out(
        n3007) );
  nor2 U2886 ( .a(n865), .b(\mat_kron/mult_40_G2_G1_G2_G2/ab[3][3] ), .out(
        n3008) );
  inv U2887 ( .in(n2276), .out(n874) );
  nor2 U2888 ( .a(n874), .b(\mat_kron/mult_40_G2_G1_G2_G2/ab[4][2] ), .out(
        n3009) );
  inv U2889 ( .in(n883), .out(n3010) );
  oai22 U2890 ( .a(n3010), .b(n2284), .c(n882), .d(n1702), .out(n3011) );
  nor2 U2891 ( .a(n2765), .b(\mat_kron/mult_40_G2_G1_G2_G2/ab[6][0] ), .out(
        n897) );
  xor2 U2892 ( .a(n3012), .b(n863), .out(n872) );
  xor2 U2893 ( .a(n3013), .b(n1700), .out(n2288) );
  xor2 U2894 ( .a(n3014), .b(n1697), .out(n1709) );
  xor2 U2895 ( .a(n3015), .b(n1702), .out(n896) );
  xor2 U2896 ( .a(n861), .b(n2275), .out(n1698) );
  xor2 U2897 ( .a(n859), .b(\mat_kron/mult_40_G2_G1_G2_G2/ab[2][4] ), .out(
        n1693) );
  xor2 U2898 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[3][3] ), .b(n865), .out(
        n3012) );
  xor2 U2899 ( .a(n2272), .b(\mat_kron/mult_40_G2_G1_G2_G2/ab[2][2] ), .out(
        n1701) );
  xor2 U2900 ( .a(n869), .b(n2277), .out(n3014) );
  xor2 U2901 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[4][2] ), .b(n2276), .out(
        n1703) );
  xor2 U2902 ( .a(n877), .b(n876), .out(n1706) );
  xor2 U2903 ( .a(n2281), .b(n879), .out(n3016) );
  xor2 U2904 ( .a(n2282), .b(n881), .out(n1708) );
  xor2 U2905 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[5][1] ), .b(n883), .out(
        n3015) );
  xor2 U2906 ( .a(n3011), .b(n895), .out(n3017) );
  xor2 U2907 ( .a(n3017), .b(n2592), .out(n1710) );
  xor2 U2908 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[5][0] ), .b(n894), .out(
        n1712) );
  xor2 U2909 ( .a(\mat_kron/mult_40_G2_G1_G2_G2/ab[3][0] ), .b(n2286), .out(
        n1713) );
  nor2 U2910 ( .a(n903), .b(\mat_kron/mult_40_G2_G1_G2_G1/ab[2][4] ), .out(
        n3018) );
  nor2 U2911 ( .a(n909), .b(\mat_kron/mult_40_G2_G1_G2_G1/ab[3][3] ), .out(
        n3019) );
  inv U2912 ( .in(n2294), .out(n918) );
  nor2 U2913 ( .a(n918), .b(\mat_kron/mult_40_G2_G1_G2_G1/ab[4][2] ), .out(
        n3020) );
  inv U2914 ( .in(n927), .out(n3021) );
  oai22 U2915 ( .a(n3021), .b(n2302), .c(n926), .d(n1723), .out(n3022) );
  nor2 U2916 ( .a(n2772), .b(\mat_kron/mult_40_G2_G1_G2_G1/ab[6][0] ), .out(
        n941) );
  xor2 U2917 ( .a(n3023), .b(n907), .out(n916) );
  xor2 U2918 ( .a(n3024), .b(n1721), .out(n2306) );
  xor2 U2919 ( .a(n3025), .b(n1718), .out(n1730) );
  xor2 U2920 ( .a(n3026), .b(n1723), .out(n940) );
  xor2 U2921 ( .a(n905), .b(n2293), .out(n1719) );
  xor2 U2922 ( .a(n903), .b(\mat_kron/mult_40_G2_G1_G2_G1/ab[2][4] ), .out(
        n1714) );
  xor2 U2923 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[3][3] ), .b(n909), .out(
        n3023) );
  xor2 U2924 ( .a(n2290), .b(\mat_kron/mult_40_G2_G1_G2_G1/ab[2][2] ), .out(
        n1722) );
  xor2 U2925 ( .a(n913), .b(n2295), .out(n3025) );
  xor2 U2926 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[4][2] ), .b(n2294), .out(
        n1724) );
  xor2 U2927 ( .a(n921), .b(n920), .out(n1727) );
  xor2 U2928 ( .a(n2299), .b(n923), .out(n3027) );
  xor2 U2929 ( .a(n2300), .b(n925), .out(n1729) );
  xor2 U2930 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[5][1] ), .b(n927), .out(
        n3026) );
  xor2 U2931 ( .a(n3022), .b(n939), .out(n3028) );
  xor2 U2932 ( .a(n3028), .b(n2598), .out(n1731) );
  xor2 U2933 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[5][0] ), .b(n938), .out(
        n1733) );
  xor2 U2934 ( .a(\mat_kron/mult_40_G2_G1_G2_G1/ab[3][0] ), .b(n2304), .out(
        n1734) );
  nor2 U2935 ( .a(n947), .b(\mat_kron/mult_40_G2_G1_G2/ab[2][4] ), .out(n3029)
         );
  nor2 U2936 ( .a(n953), .b(\mat_kron/mult_40_G2_G1_G2/ab[3][3] ), .out(n3030)
         );
  inv U2937 ( .in(n2312), .out(n962) );
  nor2 U2938 ( .a(n962), .b(\mat_kron/mult_40_G2_G1_G2/ab[4][2] ), .out(n3031)
         );
  inv U2939 ( .in(n971), .out(n3032) );
  oai22 U2940 ( .a(n3032), .b(n2320), .c(n970), .d(n1744), .out(n3033) );
  nor2 U2941 ( .a(n2779), .b(\mat_kron/mult_40_G2_G1_G2/ab[6][0] ), .out(n985)
         );
  xor2 U2942 ( .a(n3034), .b(n951), .out(n960) );
  xor2 U2943 ( .a(n3035), .b(n1742), .out(n2324) );
  xor2 U2944 ( .a(n3036), .b(n1739), .out(n1751) );
  xor2 U2945 ( .a(n3037), .b(n1744), .out(n984) );
  xor2 U2946 ( .a(n949), .b(n2311), .out(n1740) );
  xor2 U2947 ( .a(n947), .b(\mat_kron/mult_40_G2_G1_G2/ab[2][4] ), .out(n1735)
         );
  xor2 U2948 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[3][3] ), .b(n953), .out(n3034)
         );
  xor2 U2949 ( .a(n2308), .b(\mat_kron/mult_40_G2_G1_G2/ab[2][2] ), .out(n1743) );
  xor2 U2950 ( .a(n957), .b(n2313), .out(n3036) );
  xor2 U2951 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[4][2] ), .b(n2312), .out(n1745) );
  xor2 U2952 ( .a(n965), .b(n964), .out(n1748) );
  xor2 U2953 ( .a(n2317), .b(n967), .out(n3038) );
  xor2 U2954 ( .a(n2318), .b(n969), .out(n1750) );
  xor2 U2955 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[5][1] ), .b(n971), .out(n3037)
         );
  xor2 U2956 ( .a(n3033), .b(n983), .out(n3039) );
  xor2 U2957 ( .a(n3039), .b(n2604), .out(n1752) );
  xor2 U2958 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[5][0] ), .b(n982), .out(n1754)
         );
  xor2 U2959 ( .a(\mat_kron/mult_40_G2_G1_G2/ab[3][0] ), .b(n2322), .out(n1755) );
  nor2 U2960 ( .a(n991), .b(\mat_kron/mult_40_G2_G1_G1_G2/ab[2][4] ), .out(
        n3040) );
  nor2 U2961 ( .a(n997), .b(\mat_kron/mult_40_G2_G1_G1_G2/ab[3][3] ), .out(
        n3041) );
  inv U2962 ( .in(n2330), .out(n1006) );
  nor2 U2963 ( .a(n1006), .b(\mat_kron/mult_40_G2_G1_G1_G2/ab[4][2] ), .out(
        n3042) );
  inv U2964 ( .in(n1015), .out(n3043) );
  oai22 U2965 ( .a(n3043), .b(n2338), .c(n1014), .d(n1765), .out(n3044) );
  nor2 U2966 ( .a(n2786), .b(\mat_kron/mult_40_G2_G1_G1_G2/ab[6][0] ), .out(
        n1029) );
  xor2 U2967 ( .a(n3045), .b(n995), .out(n1004) );
  xor2 U2968 ( .a(n3046), .b(n1763), .out(n2342) );
  xor2 U2969 ( .a(n3047), .b(n1760), .out(n1772) );
  xor2 U2970 ( .a(n3048), .b(n1765), .out(n1028) );
  xor2 U2971 ( .a(n993), .b(n2329), .out(n1761) );
  xor2 U2972 ( .a(n991), .b(\mat_kron/mult_40_G2_G1_G1_G2/ab[2][4] ), .out(
        n1756) );
  xor2 U2973 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[3][3] ), .b(n997), .out(
        n3045) );
  xor2 U2974 ( .a(n2326), .b(\mat_kron/mult_40_G2_G1_G1_G2/ab[2][2] ), .out(
        n1764) );
  xor2 U2975 ( .a(n1001), .b(n2331), .out(n3047) );
  xor2 U2976 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[4][2] ), .b(n2330), .out(
        n1766) );
  xor2 U2977 ( .a(n1009), .b(n1008), .out(n1769) );
  xor2 U2978 ( .a(n2335), .b(n1011), .out(n3049) );
  xor2 U2979 ( .a(n2336), .b(n1013), .out(n1771) );
  xor2 U2980 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[5][1] ), .b(n1015), .out(
        n3048) );
  xor2 U2981 ( .a(n3044), .b(n1027), .out(n3050) );
  xor2 U2982 ( .a(n3050), .b(n2610), .out(n1773) );
  xor2 U2983 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[5][0] ), .b(n1026), .out(
        n1775) );
  xor2 U2984 ( .a(\mat_kron/mult_40_G2_G1_G1_G2/ab[3][0] ), .b(n2340), .out(
        n1776) );
  nor2 U2985 ( .a(n1035), .b(\mat_kron/mult_40_G2_G1_G1_G1/ab[2][4] ), .out(
        n3051) );
  nor2 U2986 ( .a(n1041), .b(\mat_kron/mult_40_G2_G1_G1_G1/ab[3][3] ), .out(
        n3052) );
  inv U2987 ( .in(n2348), .out(n1050) );
  nor2 U2988 ( .a(n1050), .b(\mat_kron/mult_40_G2_G1_G1_G1/ab[4][2] ), .out(
        n3053) );
  inv U2989 ( .in(n1059), .out(n3054) );
  oai22 U2990 ( .a(n3054), .b(n2356), .c(n1058), .d(n1786), .out(n3055) );
  nor2 U2991 ( .a(n2793), .b(\mat_kron/mult_40_G2_G1_G1_G1/ab[6][0] ), .out(
        n1073) );
  xor2 U2992 ( .a(n3056), .b(n1039), .out(n1048) );
  xor2 U2993 ( .a(n3057), .b(n1784), .out(n2360) );
  xor2 U2994 ( .a(n3058), .b(n1781), .out(n1793) );
  xor2 U2995 ( .a(n3059), .b(n1786), .out(n1072) );
  xor2 U2996 ( .a(n1037), .b(n2347), .out(n1782) );
  xor2 U2997 ( .a(n1035), .b(\mat_kron/mult_40_G2_G1_G1_G1/ab[2][4] ), .out(
        n1777) );
  xor2 U2998 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[3][3] ), .b(n1041), .out(
        n3056) );
  xor2 U2999 ( .a(n2344), .b(\mat_kron/mult_40_G2_G1_G1_G1/ab[2][2] ), .out(
        n1785) );
  xor2 U3000 ( .a(n1045), .b(n2349), .out(n3058) );
  xor2 U3001 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[4][2] ), .b(n2348), .out(
        n1787) );
  xor2 U3002 ( .a(n1053), .b(n1052), .out(n1790) );
  xor2 U3003 ( .a(n2353), .b(n1055), .out(n3060) );
  xor2 U3004 ( .a(n2354), .b(n1057), .out(n1792) );
  xor2 U3005 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[5][1] ), .b(n1059), .out(
        n3059) );
  xor2 U3006 ( .a(n3055), .b(n1071), .out(n3061) );
  xor2 U3007 ( .a(n3061), .b(n2616), .out(n1794) );
  xor2 U3008 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[5][0] ), .b(n1070), .out(
        n1796) );
  xor2 U3009 ( .a(\mat_kron/mult_40_G2_G1_G1_G1/ab[3][0] ), .b(n2358), .out(
        n1797) );
  nor2 U3010 ( .a(n1079), .b(\mat_kron/mult_40_G2_G1_G1/ab[2][4] ), .out(n3062) );
  nor2 U3011 ( .a(n1085), .b(\mat_kron/mult_40_G2_G1_G1/ab[3][3] ), .out(n3063) );
  inv U3012 ( .in(n2366), .out(n1094) );
  nor2 U3013 ( .a(n1094), .b(\mat_kron/mult_40_G2_G1_G1/ab[4][2] ), .out(n3064) );
  inv U3014 ( .in(n1103), .out(n3065) );
  oai22 U3015 ( .a(n3065), .b(n2374), .c(n1102), .d(n1807), .out(n3066) );
  nor2 U3016 ( .a(n2800), .b(\mat_kron/mult_40_G2_G1_G1/ab[6][0] ), .out(n1117) );
  xor2 U3017 ( .a(n3067), .b(n1083), .out(n1092) );
  xor2 U3018 ( .a(n3068), .b(n1805), .out(n2378) );
  xor2 U3019 ( .a(n3069), .b(n1802), .out(n1814) );
  xor2 U3020 ( .a(n3070), .b(n1807), .out(n1116) );
  xor2 U3021 ( .a(n1081), .b(n2365), .out(n1803) );
  xor2 U3022 ( .a(n1079), .b(\mat_kron/mult_40_G2_G1_G1/ab[2][4] ), .out(n1798) );
  xor2 U3023 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[3][3] ), .b(n1085), .out(n3067) );
  xor2 U3024 ( .a(n2362), .b(\mat_kron/mult_40_G2_G1_G1/ab[2][2] ), .out(n1806) );
  xor2 U3025 ( .a(n1089), .b(n2367), .out(n3069) );
  xor2 U3026 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[4][2] ), .b(n2366), .out(n1808) );
  xor2 U3027 ( .a(n1097), .b(n1096), .out(n1811) );
  xor2 U3028 ( .a(n2371), .b(n1099), .out(n3071) );
  xor2 U3029 ( .a(n2372), .b(n1101), .out(n1813) );
  xor2 U3030 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[5][1] ), .b(n1103), .out(n3070) );
  xor2 U3031 ( .a(n3066), .b(n1115), .out(n3072) );
  xor2 U3032 ( .a(n3072), .b(n2622), .out(n1815) );
  xor2 U3033 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[5][0] ), .b(n1114), .out(n1817) );
  xor2 U3034 ( .a(\mat_kron/mult_40_G2_G1_G1/ab[3][0] ), .b(n2376), .out(n1818) );
  nor2 U3035 ( .a(n1123), .b(\mat_kron/mult_40_G2_G1/ab[2][4] ), .out(n3073)
         );
  nor2 U3036 ( .a(n1129), .b(\mat_kron/mult_40_G2_G1/ab[3][3] ), .out(n3074)
         );
  inv U3037 ( .in(n2384), .out(n1138) );
  nor2 U3038 ( .a(n1138), .b(\mat_kron/mult_40_G2_G1/ab[4][2] ), .out(n3075)
         );
  inv U3039 ( .in(n1147), .out(n3076) );
  oai22 U3040 ( .a(n3076), .b(n2392), .c(n1146), .d(n1828), .out(n3077) );
  nor2 U3041 ( .a(n2807), .b(\mat_kron/mult_40_G2_G1/ab[6][0] ), .out(n1161)
         );
  xor2 U3042 ( .a(n3078), .b(n1127), .out(n1136) );
  xor2 U3043 ( .a(n3079), .b(n1826), .out(n2396) );
  xor2 U3044 ( .a(n3080), .b(n1823), .out(n1835) );
  xor2 U3045 ( .a(n3081), .b(n1828), .out(n1160) );
  xor2 U3046 ( .a(n1125), .b(n2383), .out(n1824) );
  xor2 U3047 ( .a(n1123), .b(\mat_kron/mult_40_G2_G1/ab[2][4] ), .out(n1819)
         );
  xor2 U3048 ( .a(\mat_kron/mult_40_G2_G1/ab[3][3] ), .b(n1129), .out(n3078)
         );
  xor2 U3049 ( .a(n2380), .b(\mat_kron/mult_40_G2_G1/ab[2][2] ), .out(n1827)
         );
  xor2 U3050 ( .a(n1133), .b(n2385), .out(n3080) );
  xor2 U3051 ( .a(\mat_kron/mult_40_G2_G1/ab[4][2] ), .b(n2384), .out(n1829)
         );
  xor2 U3052 ( .a(n1141), .b(n1140), .out(n1832) );
  xor2 U3053 ( .a(n2389), .b(n1143), .out(n3082) );
  xor2 U3054 ( .a(n2390), .b(n1145), .out(n1834) );
  xor2 U3055 ( .a(\mat_kron/mult_40_G2_G1/ab[5][1] ), .b(n1147), .out(n3081)
         );
  xor2 U3056 ( .a(n3077), .b(n1159), .out(n3083) );
  xor2 U3057 ( .a(n3083), .b(n2628), .out(n1836) );
  xor2 U3058 ( .a(\mat_kron/mult_40_G2_G1/ab[5][0] ), .b(n1158), .out(n1838)
         );
  xor2 U3059 ( .a(\mat_kron/mult_40_G2_G1/ab[3][0] ), .b(n2394), .out(n1839)
         );
  nor2 U3060 ( .a(n1167), .b(\mat_kron/mult_40_G2/ab[2][4] ), .out(n3084) );
  nor2 U3061 ( .a(n1173), .b(\mat_kron/mult_40_G2/ab[3][3] ), .out(n3085) );
  inv U3062 ( .in(n2402), .out(n1182) );
  nor2 U3063 ( .a(n1182), .b(\mat_kron/mult_40_G2/ab[4][2] ), .out(n3086) );
  inv U3064 ( .in(n1191), .out(n3087) );
  oai22 U3065 ( .a(n3087), .b(n2410), .c(n1190), .d(n1849), .out(n3088) );
  nor2 U3066 ( .a(n2814), .b(\mat_kron/mult_40_G2/ab[6][0] ), .out(n1205) );
  xor2 U3067 ( .a(n3089), .b(n1171), .out(n1180) );
  xor2 U3068 ( .a(n3090), .b(n1847), .out(n2414) );
  xor2 U3069 ( .a(n3091), .b(n1844), .out(n1856) );
  xor2 U3070 ( .a(n3092), .b(n1849), .out(n1204) );
  xor2 U3071 ( .a(n1169), .b(n2401), .out(n1845) );
  xor2 U3072 ( .a(n1167), .b(\mat_kron/mult_40_G2/ab[2][4] ), .out(n1840) );
  xor2 U3073 ( .a(\mat_kron/mult_40_G2/ab[3][3] ), .b(n1173), .out(n3089) );
  xor2 U3074 ( .a(n2398), .b(\mat_kron/mult_40_G2/ab[2][2] ), .out(n1848) );
  xor2 U3075 ( .a(n1177), .b(n2403), .out(n3091) );
  xor2 U3076 ( .a(\mat_kron/mult_40_G2/ab[4][2] ), .b(n2402), .out(n1850) );
  xor2 U3077 ( .a(n1185), .b(n1184), .out(n1853) );
  xor2 U3078 ( .a(n2407), .b(n1187), .out(n3093) );
  xor2 U3079 ( .a(n2408), .b(n1189), .out(n1855) );
  xor2 U3080 ( .a(\mat_kron/mult_40_G2/ab[5][1] ), .b(n1191), .out(n3092) );
  xor2 U3081 ( .a(n3088), .b(n1203), .out(n3094) );
  xor2 U3082 ( .a(n3094), .b(n2634), .out(n1857) );
  xor2 U3083 ( .a(\mat_kron/mult_40_G2/ab[5][0] ), .b(n1202), .out(n1859) );
  xor2 U3084 ( .a(\mat_kron/mult_40_G2/ab[3][0] ), .b(n2412), .out(n1860) );
  nor2 U3085 ( .a(n1211), .b(\mat_kron/mult_40/ab[2][4] ), .out(n3095) );
  nor2 U3086 ( .a(n1217), .b(\mat_kron/mult_40/ab[3][3] ), .out(n3096) );
  inv U3087 ( .in(n2420), .out(n1226) );
  nor2 U3088 ( .a(n1226), .b(\mat_kron/mult_40/ab[4][2] ), .out(n3097) );
  inv U3089 ( .in(n1235), .out(n3098) );
  oai22 U3090 ( .a(n3098), .b(n2428), .c(n1234), .d(n1870), .out(n3099) );
  nor2 U3091 ( .a(n2821), .b(\mat_kron/mult_40/ab[6][0] ), .out(n1249) );
  xor2 U3092 ( .a(n3100), .b(n1215), .out(n1224) );
  xor2 U3093 ( .a(n3101), .b(n1868), .out(n2432) );
  xor2 U3094 ( .a(n3102), .b(n1865), .out(n1877) );
  xor2 U3095 ( .a(n3103), .b(n1870), .out(n1248) );
  xor2 U3096 ( .a(n1213), .b(n2419), .out(n1866) );
  xor2 U3097 ( .a(n1211), .b(\mat_kron/mult_40/ab[2][4] ), .out(n1861) );
  xor2 U3098 ( .a(\mat_kron/mult_40/ab[3][3] ), .b(n1217), .out(n3100) );
  xor2 U3099 ( .a(n2416), .b(\mat_kron/mult_40/ab[2][2] ), .out(n1869) );
  xor2 U3100 ( .a(n1221), .b(n2421), .out(n3102) );
  xor2 U3101 ( .a(\mat_kron/mult_40/ab[4][2] ), .b(n2420), .out(n1871) );
  xor2 U3102 ( .a(n1229), .b(n1228), .out(n1874) );
  xor2 U3103 ( .a(n2425), .b(n1231), .out(n3104) );
  xor2 U3104 ( .a(n2426), .b(n1233), .out(n1876) );
  xor2 U3105 ( .a(\mat_kron/mult_40/ab[5][1] ), .b(n1235), .out(n3103) );
  xor2 U3106 ( .a(n3099), .b(n1247), .out(n3105) );
  xor2 U3107 ( .a(n3105), .b(n2640), .out(n1878) );
  xor2 U3108 ( .a(\mat_kron/mult_40/ab[5][0] ), .b(n1246), .out(n1880) );
  xor2 U3109 ( .a(\mat_kron/mult_40/ab[3][0] ), .b(n2430), .out(n1881) );
  inv U3110 ( .in(A[15]), .out(n3106) );
  inv U3111 ( .in(n191), .out(n1298) );
  nor2 U3112 ( .a(n1313), .b(\mat_sub/r102/B_AS [6]), .out(n3107) );
  oai22 U3113 ( .a(n2434), .b(n2487), .c(n1370), .d(n2486), .out(n2000) );
  aoi22 U3114 ( .a(A[10]), .b(\mat_add/r102/B_AS [2]), .c(n2000), .d(n3108), 
        .out(n1999) );
  oai22 U3115 ( .a(n2461), .b(n2500), .c(n1999), .d(n1372), .out(n1996) );
  aoi22 U3116 ( .a(A[12]), .b(\mat_add/r102/B_AS [4]), .c(n1996), .d(n3109), 
        .out(n1995) );
  oai22 U3117 ( .a(n2464), .b(n2501), .c(n1995), .d(n1374), .out(n1377) );
  nor2 U3118 ( .a(A[14]), .b(\mat_add/r102/B_AS [6]), .out(n3110) );
  xor2 U3119 ( .a(n3106), .b(\mat_sub/r102/B_AS [7]), .out(n1904) );
  xor2 U3120 ( .a(\mat_sub/r102/B_AS [6]), .b(A[14]), .out(n1905) );
  xor2 U3121 ( .a(\mat_sub/r102/B_AS [5]), .b(n2464), .out(n1906) );
  xor2 U3122 ( .a(n1306), .b(A[12]), .out(n1907) );
  xor2 U3123 ( .a(n1303), .b(A[11]), .out(n1908) );
  xor2 U3124 ( .a(n1300), .b(A[10]), .out(n1909) );
  xor2 U3125 ( .a(n2486), .b(A[9]), .out(n2650) );
  xor2 U3126 ( .a(n3106), .b(\mat_add/r102/B_AS [7]), .out(n1992) );
  xor2 U3127 ( .a(\mat_add/r102/B_AS [5]), .b(n2464), .out(n1994) );
  xor2 U3128 ( .a(\mat_add/r102/B_AS [3]), .b(n2461), .out(n1998) );
  inv U3129 ( .in(A[7]), .out(n3111) );
  inv U3130 ( .in(n195), .out(n1253) );
  nor2 U3131 ( .a(n1266), .b(\mat_sub/r106/B_AS [6]), .out(n3112) );
  oai22 U3132 ( .a(n2435), .b(n2489), .c(n1346), .d(n2488), .out(n1972) );
  aoi22 U3133 ( .a(A[2]), .b(\mat_add/r106/B_AS [2]), .c(n1972), .d(n3113), 
        .out(n1969) );
  oai22 U3134 ( .a(n2438), .b(n2490), .c(n1969), .d(n1348), .out(n1966) );
  aoi22 U3135 ( .a(A[4]), .b(\mat_add/r106/B_AS [4]), .c(n1966), .d(n3114), 
        .out(n1965) );
  oai22 U3136 ( .a(n2441), .b(n2491), .c(n1965), .d(n1350), .out(n1353) );
  nor2 U3137 ( .a(A[6]), .b(\mat_add/r106/B_AS [6]), .out(n3115) );
  xor2 U3138 ( .a(n3111), .b(\mat_sub/r106/B_AS [7]), .out(n1883) );
  xor2 U3139 ( .a(\mat_sub/r106/B_AS [6]), .b(A[6]), .out(n1884) );
  xor2 U3140 ( .a(\mat_sub/r106/B_AS [5]), .b(n2441), .out(n1885) );
  xor2 U3141 ( .a(\mat_sub/r106/B_AS [4]), .b(A[4]), .out(n1886) );
  xor2 U3142 ( .a(\mat_sub/r106/B_AS [3]), .b(n2438), .out(n1887) );
  xor2 U3143 ( .a(\mat_sub/r106/B_AS [2]), .b(A[2]), .out(n1890) );
  xor2 U3144 ( .a(n3111), .b(\mat_add/r106/B_AS [7]), .out(n1962) );
  xor2 U3145 ( .a(\mat_add/r106/B_AS [5]), .b(n2441), .out(n1964) );
  xor2 U3146 ( .a(\mat_add/r106/B_AS [3]), .b(n2438), .out(n1968) );
  xor2 U3147 ( .a(n2488), .b(A[1]), .out(n2652) );
  inv U3148 ( .in(A[31]), .out(n3116) );
  inv U3149 ( .in(n193), .out(n1268) );
  nor2 U3150 ( .a(n1281), .b(\mat_sub/r94/B_AS [6]), .out(n3117) );
  oai22 U3151 ( .a(n2443), .b(n2493), .c(n1354), .d(n2492), .out(n1980) );
  aoi22 U3152 ( .a(A[26]), .b(\mat_add/r94/B_AS [2]), .c(n1980), .d(n3118), 
        .out(n1979) );
  oai22 U3153 ( .a(n2446), .b(n2494), .c(n1979), .d(n1356), .out(n1976) );
  aoi22 U3154 ( .a(A[28]), .b(\mat_add/r94/B_AS [4]), .c(n1976), .d(n3119), 
        .out(n1975) );
  oai22 U3155 ( .a(n2449), .b(n2495), .c(n1975), .d(n1358), .out(n1361) );
  nor2 U3156 ( .a(A[30]), .b(\mat_add/r94/B_AS [6]), .out(n3120) );
  xor2 U3157 ( .a(n3116), .b(\mat_sub/r94/B_AS [7]), .out(n1888) );
  xor2 U3158 ( .a(\mat_sub/r94/B_AS [6]), .b(A[30]), .out(n1889) );
  xor2 U3159 ( .a(\mat_sub/r94/B_AS [5]), .b(n2449), .out(n1891) );
  xor2 U3160 ( .a(\mat_sub/r94/B_AS [4]), .b(A[28]), .out(n1892) );
  xor2 U3161 ( .a(\mat_sub/r94/B_AS [3]), .b(n2446), .out(n1893) );
  xor2 U3162 ( .a(\mat_sub/r94/B_AS [2]), .b(A[26]), .out(n1894) );
  xor2 U3163 ( .a(n3116), .b(\mat_add/r94/B_AS [7]), .out(n1970) );
  xor2 U3164 ( .a(\mat_add/r94/B_AS [5]), .b(n2449), .out(n1974) );
  xor2 U3165 ( .a(\mat_add/r94/B_AS [3]), .b(n2446), .out(n1978) );
  xor2 U3166 ( .a(n2492), .b(A[25]), .out(n2651) );
  inv U3167 ( .in(A[23]), .out(n3121) );
  inv U3168 ( .in(n189), .out(n1283) );
  nor2 U3169 ( .a(n1296), .b(\mat_sub/r98/B_AS [6]), .out(n3122) );
  oai22 U3170 ( .a(n2451), .b(n2497), .c(n1362), .d(n2496), .out(n1990) );
  aoi22 U3171 ( .a(A[18]), .b(\mat_add/r98/B_AS [2]), .c(n1990), .d(n3123), 
        .out(n1989) );
  oai22 U3172 ( .a(n2454), .b(n2498), .c(n1989), .d(n1364), .out(n1986) );
  aoi22 U3173 ( .a(A[20]), .b(\mat_add/r98/B_AS [4]), .c(n1986), .d(n3124), 
        .out(n1985) );
  oai22 U3174 ( .a(n2457), .b(n2499), .c(n1985), .d(n1366), .out(n1369) );
  nor2 U3175 ( .a(A[22]), .b(\mat_add/r98/B_AS [6]), .out(n3125) );
  xor2 U3176 ( .a(n3121), .b(\mat_sub/r98/B_AS [7]), .out(n1896) );
  xor2 U3177 ( .a(\mat_sub/r98/B_AS [6]), .b(A[22]), .out(n1897) );
  xor2 U3178 ( .a(\mat_sub/r98/B_AS [5]), .b(n2457), .out(n1898) );
  xor2 U3179 ( .a(\mat_sub/r98/B_AS [4]), .b(A[20]), .out(n1899) );
  xor2 U3180 ( .a(\mat_sub/r98/B_AS [3]), .b(n2454), .out(n1901) );
  xor2 U3181 ( .a(\mat_sub/r98/B_AS [2]), .b(A[18]), .out(n1902) );
  xor2 U3182 ( .a(n3121), .b(\mat_add/r98/B_AS [7]), .out(n1982) );
  xor2 U3183 ( .a(\mat_add/r98/B_AS [5]), .b(n2457), .out(n1984) );
  xor2 U3184 ( .a(\mat_add/r98/B_AS [3]), .b(n2454), .out(n1988) );
  xor2 U3185 ( .a(n2496), .b(A[17]), .out(n2653) );
  inv U3186 ( .in(n217), .out(n2010) );
  inv U3187 ( .in(n226), .out(n2015) );
  inv U3188 ( .in(n229), .out(n2016) );
  inv U3189 ( .in(\mat_mul/mult_37_G2_G2_G2/ab[6][0] ), .out(n238) );
  inv U3190 ( .in(n2827), .out(n204) );
  inv U3191 ( .in(n261), .out(n2028) );
  inv U3192 ( .in(n270), .out(n2033) );
  inv U3193 ( .in(n273), .out(n2034) );
  inv U3194 ( .in(\mat_mul/mult_37_G2_G2_G1/ab[6][0] ), .out(n282) );
  inv U3195 ( .in(n2853), .out(n248) );
  inv U3196 ( .in(n305), .out(n2046) );
  inv U3197 ( .in(n314), .out(n2051) );
  inv U3198 ( .in(n317), .out(n2052) );
  inv U3199 ( .in(\mat_mul/mult_37_G2_G2/ab[6][0] ), .out(n326) );
  inv U3200 ( .in(n2832), .out(n292) );
  inv U3201 ( .in(n349), .out(n2064) );
  inv U3202 ( .in(n358), .out(n2069) );
  inv U3203 ( .in(n361), .out(n2070) );
  inv U3204 ( .in(\mat_mul/mult_37_G2_G1_G2/ab[6][0] ), .out(n370) );
  inv U3205 ( .in(n2879), .out(n336) );
  inv U3206 ( .in(n393), .out(n2082) );
  inv U3207 ( .in(n402), .out(n2087) );
  inv U3208 ( .in(n405), .out(n2088) );
  inv U3209 ( .in(\mat_mul/mult_37_G2_G1_G1/ab[6][0] ), .out(n414) );
  inv U3210 ( .in(n2905), .out(n380) );
  inv U3211 ( .in(n437), .out(n2100) );
  inv U3212 ( .in(n446), .out(n2105) );
  inv U3213 ( .in(n449), .out(n2106) );
  inv U3214 ( .in(\mat_mul/mult_37_G2_G1/ab[6][0] ), .out(n458) );
  inv U3215 ( .in(n2858), .out(n424) );
  inv U3216 ( .in(n481), .out(n2118) );
  inv U3217 ( .in(n490), .out(n2123) );
  inv U3218 ( .in(n493), .out(n2124) );
  inv U3219 ( .in(\mat_mul/mult_37_G2/ab[6][0] ), .out(n502) );
  inv U3220 ( .in(n2884), .out(n468) );
  inv U3221 ( .in(n525), .out(n2136) );
  inv U3222 ( .in(n534), .out(n2141) );
  inv U3223 ( .in(n537), .out(n2142) );
  inv U3224 ( .in(\mat_mul/mult_37/ab[6][0] ), .out(n546) );
  inv U3225 ( .in(n2910), .out(n512) );
  inv U3226 ( .in(n569), .out(n2154) );
  inv U3227 ( .in(n578), .out(n2159) );
  inv U3228 ( .in(n581), .out(n2160) );
  inv U3229 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/ab[6][0] ), .out(n590) );
  inv U3230 ( .in(n2931), .out(n556) );
  inv U3231 ( .in(n613), .out(n2172) );
  inv U3232 ( .in(n622), .out(n2177) );
  inv U3233 ( .in(n625), .out(n2178) );
  inv U3234 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/ab[6][0] ), .out(n634) );
  inv U3235 ( .in(n2942), .out(n600) );
  inv U3236 ( .in(n657), .out(n2190) );
  inv U3237 ( .in(n666), .out(n2195) );
  inv U3238 ( .in(n669), .out(n2196) );
  inv U3239 ( .in(\mat_kron/mult_40_G2_G2_G2/ab[6][0] ), .out(n678) );
  inv U3240 ( .in(n2953), .out(n644) );
  inv U3241 ( .in(n701), .out(n2208) );
  inv U3242 ( .in(n710), .out(n2213) );
  inv U3243 ( .in(n713), .out(n2214) );
  inv U3244 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/ab[6][0] ), .out(n722) );
  inv U3245 ( .in(n2964), .out(n688) );
  inv U3246 ( .in(n745), .out(n2226) );
  inv U3247 ( .in(n754), .out(n2231) );
  inv U3248 ( .in(n757), .out(n2232) );
  inv U3249 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/ab[6][0] ), .out(n766) );
  inv U3250 ( .in(n2975), .out(n732) );
  inv U3251 ( .in(n789), .out(n2244) );
  inv U3252 ( .in(n798), .out(n2249) );
  inv U3253 ( .in(n801), .out(n2250) );
  inv U3254 ( .in(\mat_kron/mult_40_G2_G2_G1/ab[6][0] ), .out(n810) );
  inv U3255 ( .in(n2986), .out(n776) );
  inv U3256 ( .in(n833), .out(n2262) );
  inv U3257 ( .in(n842), .out(n2267) );
  inv U3258 ( .in(n845), .out(n2268) );
  inv U3259 ( .in(\mat_kron/mult_40_G2_G2/ab[6][0] ), .out(n854) );
  inv U3260 ( .in(n2997), .out(n820) );
  inv U3261 ( .in(n877), .out(n2280) );
  inv U3262 ( .in(n886), .out(n2285) );
  inv U3263 ( .in(n889), .out(n2286) );
  inv U3264 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/ab[6][0] ), .out(n898) );
  inv U3265 ( .in(n3008), .out(n864) );
  inv U3266 ( .in(n921), .out(n2298) );
  inv U3267 ( .in(n930), .out(n2303) );
  inv U3268 ( .in(n933), .out(n2304) );
  inv U3269 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/ab[6][0] ), .out(n942) );
  inv U3270 ( .in(n3019), .out(n908) );
  inv U3271 ( .in(n965), .out(n2316) );
  inv U3272 ( .in(n974), .out(n2321) );
  inv U3273 ( .in(n977), .out(n2322) );
  inv U3274 ( .in(\mat_kron/mult_40_G2_G1_G2/ab[6][0] ), .out(n986) );
  inv U3275 ( .in(n3030), .out(n952) );
  inv U3276 ( .in(n1009), .out(n2334) );
  inv U3277 ( .in(n1018), .out(n2339) );
  inv U3278 ( .in(n1021), .out(n2340) );
  inv U3279 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/ab[6][0] ), .out(n1030) );
  inv U3280 ( .in(n3041), .out(n996) );
  inv U3281 ( .in(n1053), .out(n2352) );
  inv U3282 ( .in(n1062), .out(n2357) );
  inv U3283 ( .in(n1065), .out(n2358) );
  inv U3284 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/ab[6][0] ), .out(n1074) );
  inv U3285 ( .in(n3052), .out(n1040) );
  inv U3286 ( .in(n1097), .out(n2370) );
  inv U3287 ( .in(n1106), .out(n2375) );
  inv U3288 ( .in(n1109), .out(n2376) );
  inv U3289 ( .in(\mat_kron/mult_40_G2_G1_G1/ab[6][0] ), .out(n1118) );
  inv U3290 ( .in(n3063), .out(n1084) );
  inv U3291 ( .in(n1141), .out(n2388) );
  inv U3292 ( .in(n1150), .out(n2393) );
  inv U3293 ( .in(n1153), .out(n2394) );
  inv U3294 ( .in(\mat_kron/mult_40_G2_G1/ab[6][0] ), .out(n1162) );
  inv U3295 ( .in(n3074), .out(n1128) );
  inv U3296 ( .in(n1185), .out(n2406) );
  inv U3297 ( .in(n1194), .out(n2411) );
  inv U3298 ( .in(n1197), .out(n2412) );
  inv U3299 ( .in(\mat_kron/mult_40_G2/ab[6][0] ), .out(n1206) );
  inv U3300 ( .in(n3085), .out(n1172) );
  inv U3301 ( .in(n1229), .out(n2424) );
  inv U3302 ( .in(n1238), .out(n2429) );
  inv U3303 ( .in(n1241), .out(n2430) );
  inv U3304 ( .in(\mat_kron/mult_40/ab[6][0] ), .out(n1250) );
  inv U3305 ( .in(n3096), .out(n1216) );
  inv U3306 ( .in(n190), .out(m_sub[8]) );
  inv U3307 ( .in(n192), .out(m_sub[24]) );
  inv U3308 ( .in(n188), .out(m_sub[16]) );
  inv U3309 ( .in(n194), .out(m_sub[0]) );
  inv U3310 ( .in(n1317), .out(n2837) );
  inv U3311 ( .in(n1319), .out(n2838) );
  inv U3312 ( .in(n1321), .out(n2839) );
  inv U3313 ( .in(n1325), .out(n2915) );
  inv U3314 ( .in(n1327), .out(n2916) );
  inv U3315 ( .in(n1329), .out(n2917) );
  inv U3316 ( .in(n1333), .out(n2863) );
  inv U3317 ( .in(n1335), .out(n2864) );
  inv U3318 ( .in(n1337), .out(n2865) );
  inv U3319 ( .in(n1341), .out(n2889) );
  inv U3320 ( .in(n1343), .out(n2890) );
  inv U3321 ( .in(n1345), .out(n2891) );
  inv U3322 ( .in(n3115), .out(n1352) );
  inv U3323 ( .in(n3120), .out(n1360) );
  inv U3324 ( .in(n3125), .out(n1368) );
  inv U3325 ( .in(n3110), .out(n1376) );
  inv U3326 ( .in(n1371), .out(n3108) );
  inv U3327 ( .in(n1373), .out(n3109) );
  inv U3328 ( .in(n233), .out(n2019) );
  inv U3329 ( .in(n277), .out(n2037) );
  inv U3330 ( .in(n321), .out(n2055) );
  inv U3331 ( .in(n365), .out(n2073) );
  inv U3332 ( .in(n409), .out(n2091) );
  inv U3333 ( .in(n453), .out(n2109) );
  inv U3334 ( .in(n497), .out(n2127) );
  inv U3335 ( .in(n541), .out(n2145) );
  inv U3336 ( .in(n585), .out(n2163) );
  inv U3337 ( .in(n629), .out(n2181) );
  inv U3338 ( .in(n673), .out(n2199) );
  inv U3339 ( .in(n717), .out(n2217) );
  inv U3340 ( .in(n761), .out(n2235) );
  inv U3341 ( .in(n805), .out(n2253) );
  inv U3342 ( .in(n849), .out(n2271) );
  inv U3343 ( .in(n893), .out(n2289) );
  inv U3344 ( .in(n937), .out(n2307) );
  inv U3345 ( .in(n981), .out(n2325) );
  inv U3346 ( .in(n1025), .out(n2343) );
  inv U3347 ( .in(n1069), .out(n2361) );
  inv U3348 ( .in(n1113), .out(n2379) );
  inv U3349 ( .in(n1157), .out(n2397) );
  inv U3350 ( .in(n1201), .out(n2415) );
  inv U3351 ( .in(n1245), .out(n2433) );
  inv U3352 ( .in(\mat_sub/r106/B_AS [5]), .out(n1262) );
  inv U3353 ( .in(n3112), .out(n1265) );
  inv U3354 ( .in(\mat_sub/r94/B_AS [5]), .out(n1277) );
  inv U3355 ( .in(n3117), .out(n1280) );
  inv U3356 ( .in(\mat_sub/r98/B_AS [5]), .out(n1292) );
  inv U3357 ( .in(n3122), .out(n1295) );
  inv U3358 ( .in(n1301), .out(n2460) );
  inv U3359 ( .in(n1307), .out(n2463) );
  inv U3360 ( .in(n3107), .out(n1312) );
  inv U3361 ( .in(n1316), .out(n2836) );
  inv U3362 ( .in(n1315), .out(n2824) );
  inv U3363 ( .in(n1324), .out(n2914) );
  inv U3364 ( .in(n1323), .out(n2823) );
  inv U3365 ( .in(n1332), .out(n2862) );
  inv U3366 ( .in(n1331), .out(n2825) );
  inv U3367 ( .in(n210), .out(n2007) );
  inv U3368 ( .in(n254), .out(n2025) );
  inv U3369 ( .in(n298), .out(n2043) );
  inv U3370 ( .in(n342), .out(n2061) );
  inv U3371 ( .in(n386), .out(n2079) );
  inv U3372 ( .in(n430), .out(n2097) );
  inv U3373 ( .in(n474), .out(n2115) );
  inv U3374 ( .in(n518), .out(n2133) );
  inv U3375 ( .in(n562), .out(n2151) );
  inv U3376 ( .in(n606), .out(n2169) );
  inv U3377 ( .in(n650), .out(n2187) );
  inv U3378 ( .in(n694), .out(n2205) );
  inv U3379 ( .in(n738), .out(n2223) );
  inv U3380 ( .in(n782), .out(n2241) );
  inv U3381 ( .in(n826), .out(n2259) );
  inv U3382 ( .in(n870), .out(n2277) );
  inv U3383 ( .in(n914), .out(n2295) );
  inv U3384 ( .in(n958), .out(n2313) );
  inv U3385 ( .in(n1002), .out(n2331) );
  inv U3386 ( .in(n1046), .out(n2349) );
  inv U3387 ( .in(n1090), .out(n2367) );
  inv U3388 ( .in(n1134), .out(n2385) );
  inv U3389 ( .in(n1178), .out(n2403) );
  inv U3390 ( .in(n1222), .out(n2421) );
  inv U3391 ( .in(\mat_sub/r106/B_AS [1]), .out(n2436) );
  inv U3392 ( .in(\mat_sub/r106/B_AS [3]), .out(n1257) );
  inv U3393 ( .in(n1259), .out(n2440) );
  inv U3394 ( .in(\mat_sub/r94/B_AS [1]), .out(n2444) );
  inv U3395 ( .in(\mat_sub/r94/B_AS [3]), .out(n1272) );
  inv U3396 ( .in(n1274), .out(n2448) );
  inv U3397 ( .in(\mat_sub/r98/B_AS [1]), .out(n2452) );
  inv U3398 ( .in(\mat_sub/r98/B_AS [3]), .out(n1287) );
  inv U3399 ( .in(n1289), .out(n2456) );
  inv U3400 ( .in(n1347), .out(n3113) );
  inv U3401 ( .in(n1349), .out(n3114) );
  inv U3402 ( .in(n1355), .out(n3118) );
  inv U3403 ( .in(n1357), .out(n3119) );
  inv U3404 ( .in(n1363), .out(n3123) );
  inv U3405 ( .in(n1365), .out(n3124) );
  inv U3406 ( .in(n221), .out(n2013) );
  inv U3407 ( .in(n2002), .out(n207) );
  inv U3408 ( .in(n2008), .out(n199) );
  inv U3409 ( .in(n265), .out(n2031) );
  inv U3410 ( .in(n2020), .out(n251) );
  inv U3411 ( .in(n2026), .out(n243) );
  inv U3412 ( .in(n309), .out(n2049) );
  inv U3413 ( .in(n2038), .out(n295) );
  inv U3414 ( .in(n2044), .out(n287) );
  inv U3415 ( .in(n353), .out(n2067) );
  inv U3416 ( .in(n2056), .out(n339) );
  inv U3417 ( .in(n2062), .out(n331) );
  inv U3418 ( .in(n397), .out(n2085) );
  inv U3419 ( .in(n2074), .out(n383) );
  inv U3420 ( .in(n2080), .out(n375) );
  inv U3421 ( .in(n441), .out(n2103) );
  inv U3422 ( .in(n2092), .out(n427) );
  inv U3423 ( .in(n2098), .out(n419) );
  inv U3424 ( .in(n485), .out(n2121) );
  inv U3425 ( .in(n2110), .out(n471) );
  inv U3426 ( .in(n2116), .out(n463) );
  inv U3427 ( .in(n529), .out(n2139) );
  inv U3428 ( .in(n2128), .out(n515) );
  inv U3429 ( .in(n2134), .out(n507) );
  inv U3430 ( .in(n573), .out(n2157) );
  inv U3431 ( .in(n2146), .out(n559) );
  inv U3432 ( .in(n2152), .out(n551) );
  inv U3433 ( .in(n617), .out(n2175) );
  inv U3434 ( .in(n2164), .out(n603) );
  inv U3435 ( .in(n2170), .out(n595) );
  inv U3436 ( .in(n661), .out(n2193) );
  inv U3437 ( .in(n2182), .out(n647) );
  inv U3438 ( .in(n2188), .out(n639) );
  inv U3439 ( .in(n705), .out(n2211) );
  inv U3440 ( .in(n2200), .out(n691) );
  inv U3441 ( .in(n2206), .out(n683) );
  inv U3442 ( .in(n749), .out(n2229) );
  inv U3443 ( .in(n2218), .out(n735) );
  inv U3444 ( .in(n2224), .out(n727) );
  inv U3445 ( .in(n793), .out(n2247) );
  inv U3446 ( .in(n2236), .out(n779) );
  inv U3447 ( .in(n2242), .out(n771) );
  inv U3448 ( .in(n837), .out(n2265) );
  inv U3449 ( .in(n2254), .out(n823) );
  inv U3450 ( .in(n2260), .out(n815) );
  inv U3451 ( .in(n881), .out(n2283) );
  inv U3452 ( .in(n2272), .out(n867) );
  inv U3453 ( .in(n2278), .out(n859) );
  inv U3454 ( .in(n925), .out(n2301) );
  inv U3455 ( .in(n2290), .out(n911) );
  inv U3456 ( .in(n2296), .out(n903) );
  inv U3457 ( .in(n969), .out(n2319) );
  inv U3458 ( .in(n2308), .out(n955) );
  inv U3459 ( .in(n2314), .out(n947) );
  inv U3460 ( .in(n1013), .out(n2337) );
  inv U3461 ( .in(n2326), .out(n999) );
  inv U3462 ( .in(n2332), .out(n991) );
  inv U3463 ( .in(n1057), .out(n2355) );
  inv U3464 ( .in(n2344), .out(n1043) );
  inv U3465 ( .in(n2350), .out(n1035) );
  inv U3466 ( .in(n1101), .out(n2373) );
  inv U3467 ( .in(n2362), .out(n1087) );
  inv U3468 ( .in(n2368), .out(n1079) );
  inv U3469 ( .in(n1145), .out(n2391) );
  inv U3470 ( .in(n2380), .out(n1131) );
  inv U3471 ( .in(n2386), .out(n1123) );
  inv U3472 ( .in(n1189), .out(n2409) );
  inv U3473 ( .in(n2398), .out(n1175) );
  inv U3474 ( .in(n2404), .out(n1167) );
  inv U3475 ( .in(n1233), .out(n2427) );
  inv U3476 ( .in(n2416), .out(n1219) );
  inv U3477 ( .in(n2422), .out(n1211) );
  inv U3478 ( .in(n1254), .out(n2437) );
  inv U3479 ( .in(n1269), .out(n2445) );
  inv U3480 ( .in(n1284), .out(n2453) );
  inv U3481 ( .in(\mat_sub/r102/B_AS [3]), .out(n1303) );
  inv U3482 ( .in(\mat_mul/mult_37_G2_G2_G2/ab[3][1] ), .out(n2011) );
  inv U3483 ( .in(\mat_mul/mult_37_G2_G2_G2/ab[3][2] ), .out(n209) );
  inv U3484 ( .in(n2004), .out(n201) );
  inv U3485 ( .in(\mat_mul/mult_37_G2_G2_G2/ab[2][0] ), .out(n225) );
  inv U3486 ( .in(\mat_mul/mult_37_G2_G2_G2/ab[3][0] ), .out(n228) );
  inv U3487 ( .in(\mat_mul/mult_37_G2_G2_G1/ab[3][1] ), .out(n2029) );
  inv U3488 ( .in(\mat_mul/mult_37_G2_G2_G1/ab[3][2] ), .out(n253) );
  inv U3489 ( .in(n2022), .out(n245) );
  inv U3490 ( .in(\mat_mul/mult_37_G2_G2_G1/ab[2][0] ), .out(n269) );
  inv U3491 ( .in(\mat_mul/mult_37_G2_G2_G1/ab[3][0] ), .out(n272) );
  inv U3492 ( .in(\mat_mul/mult_37_G2_G2/ab[3][1] ), .out(n2047) );
  inv U3493 ( .in(\mat_mul/mult_37_G2_G2/ab[3][2] ), .out(n297) );
  inv U3494 ( .in(n2040), .out(n289) );
  inv U3495 ( .in(\mat_mul/mult_37_G2_G2/ab[2][0] ), .out(n313) );
  inv U3496 ( .in(\mat_mul/mult_37_G2_G2/ab[3][0] ), .out(n316) );
  inv U3497 ( .in(\mat_mul/mult_37_G2_G1_G2/ab[3][1] ), .out(n2065) );
  inv U3498 ( .in(\mat_mul/mult_37_G2_G1_G2/ab[3][2] ), .out(n341) );
  inv U3499 ( .in(n2058), .out(n333) );
  inv U3500 ( .in(\mat_mul/mult_37_G2_G1_G2/ab[2][0] ), .out(n357) );
  inv U3501 ( .in(\mat_mul/mult_37_G2_G1_G2/ab[3][0] ), .out(n360) );
  inv U3502 ( .in(\mat_mul/mult_37_G2_G1_G1/ab[3][1] ), .out(n2083) );
  inv U3503 ( .in(\mat_mul/mult_37_G2_G1_G1/ab[3][2] ), .out(n385) );
  inv U3504 ( .in(n2076), .out(n377) );
  inv U3505 ( .in(\mat_mul/mult_37_G2_G1_G1/ab[2][0] ), .out(n401) );
  inv U3506 ( .in(\mat_mul/mult_37_G2_G1_G1/ab[3][0] ), .out(n404) );
  inv U3507 ( .in(\mat_mul/mult_37_G2_G1/ab[3][1] ), .out(n2101) );
  inv U3508 ( .in(\mat_mul/mult_37_G2_G1/ab[3][2] ), .out(n429) );
  inv U3509 ( .in(n2094), .out(n421) );
  inv U3510 ( .in(\mat_mul/mult_37_G2_G1/ab[2][0] ), .out(n445) );
  inv U3511 ( .in(\mat_mul/mult_37_G2_G1/ab[3][0] ), .out(n448) );
  inv U3512 ( .in(\mat_mul/mult_37_G2/ab[3][1] ), .out(n2119) );
  inv U3513 ( .in(\mat_mul/mult_37_G2/ab[3][2] ), .out(n473) );
  inv U3514 ( .in(n2112), .out(n465) );
  inv U3515 ( .in(\mat_mul/mult_37_G2/ab[2][0] ), .out(n489) );
  inv U3516 ( .in(\mat_mul/mult_37_G2/ab[3][0] ), .out(n492) );
  inv U3517 ( .in(\mat_mul/mult_37/ab[3][1] ), .out(n2137) );
  inv U3518 ( .in(\mat_mul/mult_37/ab[3][2] ), .out(n517) );
  inv U3519 ( .in(n2130), .out(n509) );
  inv U3520 ( .in(\mat_mul/mult_37/ab[2][0] ), .out(n533) );
  inv U3521 ( .in(\mat_mul/mult_37/ab[3][0] ), .out(n536) );
  inv U3522 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/ab[3][1] ), .out(n2155) );
  inv U3523 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/ab[3][2] ), .out(n561) );
  inv U3524 ( .in(n2148), .out(n553) );
  inv U3525 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/ab[2][0] ), .out(n577) );
  inv U3526 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/ab[3][0] ), .out(n580) );
  inv U3527 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/ab[3][1] ), .out(n2173) );
  inv U3528 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/ab[3][2] ), .out(n605) );
  inv U3529 ( .in(n2166), .out(n597) );
  inv U3530 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/ab[2][0] ), .out(n621) );
  inv U3531 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/ab[3][0] ), .out(n624) );
  inv U3532 ( .in(\mat_kron/mult_40_G2_G2_G2/ab[3][1] ), .out(n2191) );
  inv U3533 ( .in(\mat_kron/mult_40_G2_G2_G2/ab[3][2] ), .out(n649) );
  inv U3534 ( .in(n2184), .out(n641) );
  inv U3535 ( .in(\mat_kron/mult_40_G2_G2_G2/ab[2][0] ), .out(n665) );
  inv U3536 ( .in(\mat_kron/mult_40_G2_G2_G2/ab[3][0] ), .out(n668) );
  inv U3537 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/ab[3][1] ), .out(n2209) );
  inv U3538 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/ab[3][2] ), .out(n693) );
  inv U3539 ( .in(n2202), .out(n685) );
  inv U3540 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/ab[2][0] ), .out(n709) );
  inv U3541 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/ab[3][0] ), .out(n712) );
  inv U3542 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/ab[3][1] ), .out(n2227) );
  inv U3543 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/ab[3][2] ), .out(n737) );
  inv U3544 ( .in(n2220), .out(n729) );
  inv U3545 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/ab[2][0] ), .out(n753) );
  inv U3546 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/ab[3][0] ), .out(n756) );
  inv U3547 ( .in(\mat_kron/mult_40_G2_G2_G1/ab[3][1] ), .out(n2245) );
  inv U3548 ( .in(\mat_kron/mult_40_G2_G2_G1/ab[3][2] ), .out(n781) );
  inv U3549 ( .in(n2238), .out(n773) );
  inv U3550 ( .in(\mat_kron/mult_40_G2_G2_G1/ab[2][0] ), .out(n797) );
  inv U3551 ( .in(\mat_kron/mult_40_G2_G2_G1/ab[3][0] ), .out(n800) );
  inv U3552 ( .in(\mat_kron/mult_40_G2_G2/ab[3][1] ), .out(n2263) );
  inv U3553 ( .in(\mat_kron/mult_40_G2_G2/ab[3][2] ), .out(n825) );
  inv U3554 ( .in(n2256), .out(n817) );
  inv U3555 ( .in(\mat_kron/mult_40_G2_G2/ab[2][0] ), .out(n841) );
  inv U3556 ( .in(\mat_kron/mult_40_G2_G2/ab[3][0] ), .out(n844) );
  inv U3557 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/ab[3][1] ), .out(n2281) );
  inv U3558 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/ab[3][2] ), .out(n869) );
  inv U3559 ( .in(n2274), .out(n861) );
  inv U3560 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/ab[2][0] ), .out(n885) );
  inv U3561 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/ab[3][0] ), .out(n888) );
  inv U3562 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/ab[3][1] ), .out(n2299) );
  inv U3563 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/ab[3][2] ), .out(n913) );
  inv U3564 ( .in(n2292), .out(n905) );
  inv U3565 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/ab[2][0] ), .out(n929) );
  inv U3566 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/ab[3][0] ), .out(n932) );
  inv U3567 ( .in(\mat_kron/mult_40_G2_G1_G2/ab[3][1] ), .out(n2317) );
  inv U3568 ( .in(\mat_kron/mult_40_G2_G1_G2/ab[3][2] ), .out(n957) );
  inv U3569 ( .in(n2310), .out(n949) );
  inv U3570 ( .in(\mat_kron/mult_40_G2_G1_G2/ab[2][0] ), .out(n973) );
  inv U3571 ( .in(\mat_kron/mult_40_G2_G1_G2/ab[3][0] ), .out(n976) );
  inv U3572 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/ab[3][1] ), .out(n2335) );
  inv U3573 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/ab[3][2] ), .out(n1001) );
  inv U3574 ( .in(n2328), .out(n993) );
  inv U3575 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/ab[2][0] ), .out(n1017) );
  inv U3576 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/ab[3][0] ), .out(n1020) );
  inv U3577 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/ab[3][1] ), .out(n2353) );
  inv U3578 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/ab[3][2] ), .out(n1045) );
  inv U3579 ( .in(n2346), .out(n1037) );
  inv U3580 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/ab[2][0] ), .out(n1061) );
  inv U3581 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/ab[3][0] ), .out(n1064) );
  inv U3582 ( .in(\mat_kron/mult_40_G2_G1_G1/ab[3][1] ), .out(n2371) );
  inv U3583 ( .in(\mat_kron/mult_40_G2_G1_G1/ab[3][2] ), .out(n1089) );
  inv U3584 ( .in(n2364), .out(n1081) );
  inv U3585 ( .in(\mat_kron/mult_40_G2_G1_G1/ab[2][0] ), .out(n1105) );
  inv U3586 ( .in(\mat_kron/mult_40_G2_G1_G1/ab[3][0] ), .out(n1108) );
  inv U3587 ( .in(\mat_kron/mult_40_G2_G1/ab[3][1] ), .out(n2389) );
  inv U3588 ( .in(\mat_kron/mult_40_G2_G1/ab[3][2] ), .out(n1133) );
  inv U3589 ( .in(n2382), .out(n1125) );
  inv U3590 ( .in(\mat_kron/mult_40_G2_G1/ab[2][0] ), .out(n1149) );
  inv U3591 ( .in(\mat_kron/mult_40_G2_G1/ab[3][0] ), .out(n1152) );
  inv U3592 ( .in(\mat_kron/mult_40_G2/ab[3][1] ), .out(n2407) );
  inv U3593 ( .in(\mat_kron/mult_40_G2/ab[3][2] ), .out(n1177) );
  inv U3594 ( .in(n2400), .out(n1169) );
  inv U3595 ( .in(\mat_kron/mult_40_G2/ab[2][0] ), .out(n1193) );
  inv U3596 ( .in(\mat_kron/mult_40_G2/ab[3][0] ), .out(n1196) );
  inv U3597 ( .in(\mat_kron/mult_40/ab[3][1] ), .out(n2425) );
  inv U3598 ( .in(\mat_kron/mult_40/ab[3][2] ), .out(n1221) );
  inv U3599 ( .in(n2418), .out(n1213) );
  inv U3600 ( .in(\mat_kron/mult_40/ab[2][0] ), .out(n1237) );
  inv U3601 ( .in(\mat_kron/mult_40/ab[3][0] ), .out(n1240) );
  inv U3602 ( .in(\mat_mul/mult_37_G2_G2_G2/ab[2][1] ), .out(n216) );
  inv U3603 ( .in(n2009), .out(n219) );
  inv U3604 ( .in(n206), .out(n2003) );
  inv U3605 ( .in(\mat_mul/mult_37_G2_G2_G2/ab[1][4] ), .out(n1380) );
  inv U3606 ( .in(n230), .out(n2017) );
  inv U3607 ( .in(n2848), .out(n2841) );
  inv U3608 ( .in(n239), .out(n2660) );
  inv U3609 ( .in(n2826), .out(n198) );
  inv U3610 ( .in(n2828), .out(n213) );
  inv U3611 ( .in(\mat_mul/mult_37_G2_G2_G1/ab[2][1] ), .out(n260) );
  inv U3612 ( .in(n2027), .out(n263) );
  inv U3613 ( .in(n250), .out(n2021) );
  inv U3614 ( .in(\mat_mul/mult_37_G2_G2_G1/ab[1][4] ), .out(n1401) );
  inv U3615 ( .in(n274), .out(n2035) );
  inv U3616 ( .in(n2874), .out(n2867) );
  inv U3617 ( .in(n283), .out(n2667) );
  inv U3618 ( .in(n2852), .out(n242) );
  inv U3619 ( .in(n2854), .out(n257) );
  inv U3620 ( .in(\mat_mul/mult_37_G2_G2/ab[2][1] ), .out(n304) );
  inv U3621 ( .in(n2045), .out(n307) );
  inv U3622 ( .in(n294), .out(n2039) );
  inv U3623 ( .in(\mat_mul/mult_37_G2_G2/ab[1][4] ), .out(n1422) );
  inv U3624 ( .in(n318), .out(n2053) );
  inv U3625 ( .in(n2850), .out(n2845) );
  inv U3626 ( .in(n327), .out(n2674) );
  inv U3627 ( .in(n2831), .out(n286) );
  inv U3628 ( .in(n2833), .out(n301) );
  inv U3629 ( .in(\mat_mul/mult_37_G2_G1_G2/ab[2][1] ), .out(n348) );
  inv U3630 ( .in(n2063), .out(n351) );
  inv U3631 ( .in(n338), .out(n2057) );
  inv U3632 ( .in(\mat_mul/mult_37_G2_G1_G2/ab[1][4] ), .out(n1443) );
  inv U3633 ( .in(n362), .out(n2071) );
  inv U3634 ( .in(n2900), .out(n2893) );
  inv U3635 ( .in(n371), .out(n2681) );
  inv U3636 ( .in(n2878), .out(n330) );
  inv U3637 ( .in(n2880), .out(n345) );
  inv U3638 ( .in(\mat_mul/mult_37_G2_G1_G1/ab[2][1] ), .out(n392) );
  inv U3639 ( .in(n2081), .out(n395) );
  inv U3640 ( .in(n382), .out(n2075) );
  inv U3641 ( .in(\mat_mul/mult_37_G2_G1_G1/ab[1][4] ), .out(n1464) );
  inv U3642 ( .in(n406), .out(n2089) );
  inv U3643 ( .in(n2926), .out(n2919) );
  inv U3644 ( .in(n415), .out(n2688) );
  inv U3645 ( .in(n2904), .out(n374) );
  inv U3646 ( .in(n2906), .out(n389) );
  inv U3647 ( .in(\mat_mul/mult_37_G2_G1/ab[2][1] ), .out(n436) );
  inv U3648 ( .in(n2099), .out(n439) );
  inv U3649 ( .in(n426), .out(n2093) );
  inv U3650 ( .in(\mat_mul/mult_37_G2_G1/ab[1][4] ), .out(n1485) );
  inv U3651 ( .in(n450), .out(n2107) );
  inv U3652 ( .in(n2876), .out(n2871) );
  inv U3653 ( .in(n459), .out(n2695) );
  inv U3654 ( .in(n2857), .out(n418) );
  inv U3655 ( .in(n2859), .out(n433) );
  inv U3656 ( .in(\mat_mul/mult_37_G2/ab[2][1] ), .out(n480) );
  inv U3657 ( .in(n2117), .out(n483) );
  inv U3658 ( .in(n470), .out(n2111) );
  inv U3659 ( .in(\mat_mul/mult_37_G2/ab[1][4] ), .out(n1506) );
  inv U3660 ( .in(n494), .out(n2125) );
  inv U3661 ( .in(n2902), .out(n2897) );
  inv U3662 ( .in(n503), .out(n2702) );
  inv U3663 ( .in(n2883), .out(n462) );
  inv U3664 ( .in(n2885), .out(n477) );
  inv U3665 ( .in(\mat_mul/mult_37/ab[2][1] ), .out(n524) );
  inv U3666 ( .in(n2135), .out(n527) );
  inv U3667 ( .in(n514), .out(n2129) );
  inv U3668 ( .in(\mat_mul/mult_37/ab[1][4] ), .out(n1527) );
  inv U3669 ( .in(n538), .out(n2143) );
  inv U3670 ( .in(n2928), .out(n2923) );
  inv U3671 ( .in(n547), .out(n2709) );
  inv U3672 ( .in(n2909), .out(n506) );
  inv U3673 ( .in(n2911), .out(n521) );
  inv U3674 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/ab[2][1] ), .out(n568) );
  inv U3675 ( .in(n2153), .out(n571) );
  inv U3676 ( .in(n558), .out(n2147) );
  inv U3677 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/ab[1][4] ), .out(n1548) );
  inv U3678 ( .in(n582), .out(n2161) );
  inv U3679 ( .in(n2939), .out(n2936) );
  inv U3680 ( .in(n591), .out(n2716) );
  inv U3681 ( .in(n2930), .out(n550) );
  inv U3682 ( .in(n2932), .out(n565) );
  inv U3683 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/ab[2][1] ), .out(n612) );
  inv U3684 ( .in(n2171), .out(n615) );
  inv U3685 ( .in(n602), .out(n2165) );
  inv U3686 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/ab[1][4] ), .out(n1569) );
  inv U3687 ( .in(n626), .out(n2179) );
  inv U3688 ( .in(n2950), .out(n2947) );
  inv U3689 ( .in(n635), .out(n2723) );
  inv U3690 ( .in(n2941), .out(n594) );
  inv U3691 ( .in(n2943), .out(n609) );
  inv U3692 ( .in(\mat_kron/mult_40_G2_G2_G2/ab[2][1] ), .out(n656) );
  inv U3693 ( .in(n2189), .out(n659) );
  inv U3694 ( .in(n646), .out(n2183) );
  inv U3695 ( .in(\mat_kron/mult_40_G2_G2_G2/ab[1][4] ), .out(n1590) );
  inv U3696 ( .in(n670), .out(n2197) );
  inv U3697 ( .in(n2961), .out(n2958) );
  inv U3698 ( .in(n679), .out(n2730) );
  inv U3699 ( .in(n2952), .out(n638) );
  inv U3700 ( .in(n2954), .out(n653) );
  inv U3701 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/ab[2][1] ), .out(n700) );
  inv U3702 ( .in(n2207), .out(n703) );
  inv U3703 ( .in(n690), .out(n2201) );
  inv U3704 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/ab[1][4] ), .out(n1611) );
  inv U3705 ( .in(n714), .out(n2215) );
  inv U3706 ( .in(n2972), .out(n2969) );
  inv U3707 ( .in(n723), .out(n2737) );
  inv U3708 ( .in(n2963), .out(n682) );
  inv U3709 ( .in(n2965), .out(n697) );
  inv U3710 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/ab[2][1] ), .out(n744) );
  inv U3711 ( .in(n2225), .out(n747) );
  inv U3712 ( .in(n734), .out(n2219) );
  inv U3713 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/ab[1][4] ), .out(n1632) );
  inv U3714 ( .in(n758), .out(n2233) );
  inv U3715 ( .in(n2983), .out(n2980) );
  inv U3716 ( .in(n767), .out(n2744) );
  inv U3717 ( .in(n2974), .out(n726) );
  inv U3718 ( .in(n2976), .out(n741) );
  inv U3719 ( .in(\mat_kron/mult_40_G2_G2_G1/ab[2][1] ), .out(n788) );
  inv U3720 ( .in(n2243), .out(n791) );
  inv U3721 ( .in(n778), .out(n2237) );
  inv U3722 ( .in(\mat_kron/mult_40_G2_G2_G1/ab[1][4] ), .out(n1653) );
  inv U3723 ( .in(n802), .out(n2251) );
  inv U3724 ( .in(n2994), .out(n2991) );
  inv U3725 ( .in(n811), .out(n2751) );
  inv U3726 ( .in(n2985), .out(n770) );
  inv U3727 ( .in(n2987), .out(n785) );
  inv U3728 ( .in(\mat_kron/mult_40_G2_G2/ab[2][1] ), .out(n832) );
  inv U3729 ( .in(n2261), .out(n835) );
  inv U3730 ( .in(n822), .out(n2255) );
  inv U3731 ( .in(\mat_kron/mult_40_G2_G2/ab[1][4] ), .out(n1674) );
  inv U3732 ( .in(n846), .out(n2269) );
  inv U3733 ( .in(n3005), .out(n3002) );
  inv U3734 ( .in(n855), .out(n2758) );
  inv U3735 ( .in(n2996), .out(n814) );
  inv U3736 ( .in(n2998), .out(n829) );
  inv U3737 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/ab[2][1] ), .out(n876) );
  inv U3738 ( .in(n2279), .out(n879) );
  inv U3739 ( .in(n866), .out(n2273) );
  inv U3740 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/ab[1][4] ), .out(n1695) );
  inv U3741 ( .in(n890), .out(n2287) );
  inv U3742 ( .in(n3016), .out(n3013) );
  inv U3743 ( .in(n899), .out(n2765) );
  inv U3744 ( .in(n3007), .out(n858) );
  inv U3745 ( .in(n3009), .out(n873) );
  inv U3746 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/ab[2][1] ), .out(n920) );
  inv U3747 ( .in(n2297), .out(n923) );
  inv U3748 ( .in(n910), .out(n2291) );
  inv U3749 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/ab[1][4] ), .out(n1716) );
  inv U3750 ( .in(n934), .out(n2305) );
  inv U3751 ( .in(n3027), .out(n3024) );
  inv U3752 ( .in(n943), .out(n2772) );
  inv U3753 ( .in(n3018), .out(n902) );
  inv U3754 ( .in(n3020), .out(n917) );
  inv U3755 ( .in(\mat_kron/mult_40_G2_G1_G2/ab[2][1] ), .out(n964) );
  inv U3756 ( .in(n2315), .out(n967) );
  inv U3757 ( .in(n954), .out(n2309) );
  inv U3758 ( .in(\mat_kron/mult_40_G2_G1_G2/ab[1][4] ), .out(n1737) );
  inv U3759 ( .in(n978), .out(n2323) );
  inv U3760 ( .in(n3038), .out(n3035) );
  inv U3761 ( .in(n987), .out(n2779) );
  inv U3762 ( .in(n3029), .out(n946) );
  inv U3763 ( .in(n3031), .out(n961) );
  inv U3764 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/ab[2][1] ), .out(n1008) );
  inv U3765 ( .in(n2333), .out(n1011) );
  inv U3766 ( .in(n998), .out(n2327) );
  inv U3767 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/ab[1][4] ), .out(n1758) );
  inv U3768 ( .in(n1022), .out(n2341) );
  inv U3769 ( .in(n3049), .out(n3046) );
  inv U3770 ( .in(n1031), .out(n2786) );
  inv U3771 ( .in(n3040), .out(n990) );
  inv U3772 ( .in(n3042), .out(n1005) );
  inv U3773 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/ab[2][1] ), .out(n1052) );
  inv U3774 ( .in(n2351), .out(n1055) );
  inv U3775 ( .in(n1042), .out(n2345) );
  inv U3776 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/ab[1][4] ), .out(n1779) );
  inv U3777 ( .in(n1066), .out(n2359) );
  inv U3778 ( .in(n3060), .out(n3057) );
  inv U3779 ( .in(n1075), .out(n2793) );
  inv U3780 ( .in(n3051), .out(n1034) );
  inv U3781 ( .in(n3053), .out(n1049) );
  inv U3782 ( .in(\mat_kron/mult_40_G2_G1_G1/ab[2][1] ), .out(n1096) );
  inv U3783 ( .in(n2369), .out(n1099) );
  inv U3784 ( .in(n1086), .out(n2363) );
  inv U3785 ( .in(\mat_kron/mult_40_G2_G1_G1/ab[1][4] ), .out(n1800) );
  inv U3786 ( .in(n1110), .out(n2377) );
  inv U3787 ( .in(n3071), .out(n3068) );
  inv U3788 ( .in(n1119), .out(n2800) );
  inv U3789 ( .in(n3062), .out(n1078) );
  inv U3790 ( .in(n3064), .out(n1093) );
  inv U3791 ( .in(\mat_kron/mult_40_G2_G1/ab[2][1] ), .out(n1140) );
  inv U3792 ( .in(n2387), .out(n1143) );
  inv U3793 ( .in(n1130), .out(n2381) );
  inv U3794 ( .in(\mat_kron/mult_40_G2_G1/ab[1][4] ), .out(n1821) );
  inv U3795 ( .in(n1154), .out(n2395) );
  inv U3796 ( .in(n3082), .out(n3079) );
  inv U3797 ( .in(n1163), .out(n2807) );
  inv U3798 ( .in(n3073), .out(n1122) );
  inv U3799 ( .in(n3075), .out(n1137) );
  inv U3800 ( .in(\mat_kron/mult_40_G2/ab[2][1] ), .out(n1184) );
  inv U3801 ( .in(n2405), .out(n1187) );
  inv U3802 ( .in(n1174), .out(n2399) );
  inv U3803 ( .in(\mat_kron/mult_40_G2/ab[1][4] ), .out(n1842) );
  inv U3804 ( .in(n1198), .out(n2413) );
  inv U3805 ( .in(n3093), .out(n3090) );
  inv U3806 ( .in(n1207), .out(n2814) );
  inv U3807 ( .in(n3084), .out(n1166) );
  inv U3808 ( .in(n3086), .out(n1181) );
  inv U3809 ( .in(\mat_kron/mult_40/ab[2][1] ), .out(n1228) );
  inv U3810 ( .in(n2423), .out(n1231) );
  inv U3811 ( .in(n1218), .out(n2417) );
  inv U3812 ( .in(\mat_kron/mult_40/ab[1][4] ), .out(n1863) );
  inv U3813 ( .in(n1242), .out(n2431) );
  inv U3814 ( .in(n3104), .out(n3101) );
  inv U3815 ( .in(n1251), .out(n2821) );
  inv U3816 ( .in(n3095), .out(n1210) );
  inv U3817 ( .in(n3097), .out(n1225) );
  inv U3818 ( .in(n1256), .out(n2439) );
  inv U3819 ( .in(n1261), .out(n2442) );
  inv U3820 ( .in(n1271), .out(n2447) );
  inv U3821 ( .in(n1276), .out(n2450) );
  inv U3822 ( .in(n1286), .out(n2455) );
  inv U3823 ( .in(n1291), .out(n2458) );
  inv U3824 ( .in(n1297), .out(n2459) );
  inv U3825 ( .in(n1304), .out(n2462) );
  inv U3826 ( .in(n1308), .out(n2465) );
  inv U3827 ( .in(n1910), .out(m_mul[7]) );
  inv U3828 ( .in(n1921), .out(m_mul[31]) );
  inv U3829 ( .in(n1936), .out(m_mul[23]) );
  inv U3830 ( .in(n1949), .out(m_mul[15]) );
  inv U3831 ( .in(\mat_mul/mult_37_G2_G2_G2/A1[0] ), .out(n3126) );
  inv U3832 ( .in(n3127), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ) );
  inv U3833 ( .in(\mat_mul/mult_37_G2_G2_G2/A1[1] ), .out(n3128) );
  inv U3834 ( .in(n3129), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ) );
  inv U3835 ( .in(\mat_mul/mult_37_G2_G2_G2/A1[2] ), .out(n3130) );
  inv U3836 ( .in(n3131), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ) );
  inv U3837 ( .in(\mat_mul/mult_37_G2_G2_G2/A1[3] ), .out(n3132) );
  inv U3838 ( .in(n3133), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ) );
  inv U3839 ( .in(\mat_mul/mult_37_G2_G2_G2/A1[4] ), .out(n3134) );
  inv U3840 ( .in(n3135), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ) );
  inv U3841 ( .in(\mat_mul/mult_37_G2_G2_G2/A1[5] ), .out(n3136) );
  inv U3842 ( .in(n3137), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[7] ) );
  inv U3843 ( .in(\mat_mul/mult_37_G2_G2/A1[0] ), .out(n3138) );
  inv U3844 ( .in(n3139), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ) );
  inv U3845 ( .in(\mat_mul/mult_37_G2_G2/A1[1] ), .out(n3140) );
  inv U3846 ( .in(n3141), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[3] ) );
  inv U3847 ( .in(\mat_mul/mult_37_G2_G2/A1[2] ), .out(n3142) );
  inv U3848 ( .in(n3143), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ) );
  inv U3849 ( .in(\mat_mul/mult_37_G2_G2/A1[3] ), .out(n3144) );
  inv U3850 ( .in(n3145), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[5] ) );
  inv U3851 ( .in(\mat_mul/mult_37_G2_G2/A1[4] ), .out(n3146) );
  inv U3852 ( .in(n3147), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ) );
  inv U3853 ( .in(\mat_mul/mult_37_G2_G2/A1[5] ), .out(n3148) );
  inv U3854 ( .in(n3149), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[7] ) );
  inv U3855 ( .in(\mat_mul/mult_37_G2_G1_G2/A1[0] ), .out(n3150) );
  inv U3856 ( .in(n3151), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ) );
  inv U3857 ( .in(\mat_mul/mult_37_G2_G1_G2/A1[1] ), .out(n3152) );
  inv U3858 ( .in(n3153), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ) );
  inv U3859 ( .in(\mat_mul/mult_37_G2_G1_G2/A1[2] ), .out(n3154) );
  inv U3860 ( .in(n3155), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ) );
  inv U3861 ( .in(\mat_mul/mult_37_G2_G1_G2/A1[3] ), .out(n3156) );
  inv U3862 ( .in(n3157), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ) );
  inv U3863 ( .in(\mat_mul/mult_37_G2_G1_G2/A1[4] ), .out(n3158) );
  inv U3864 ( .in(n3159), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ) );
  inv U3865 ( .in(\mat_mul/mult_37_G2_G1_G2/A1[5] ), .out(n3160) );
  inv U3866 ( .in(n3161), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[7] ) );
  inv U3867 ( .in(\mat_mul/mult_37_G2/A1[0] ), .out(n3162) );
  inv U3868 ( .in(n3163), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ) );
  inv U3869 ( .in(\mat_mul/mult_37_G2/A1[1] ), .out(n3164) );
  inv U3870 ( .in(n3165), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[3] ) );
  inv U3871 ( .in(\mat_mul/mult_37_G2/A1[2] ), .out(n3166) );
  inv U3872 ( .in(n3167), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ) );
  inv U3873 ( .in(\mat_mul/mult_37_G2/A1[3] ), .out(n3168) );
  inv U3874 ( .in(n3169), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[5] ) );
  inv U3875 ( .in(\mat_mul/mult_37_G2/A1[4] ), .out(n3170) );
  inv U3876 ( .in(n3171), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ) );
  inv U3877 ( .in(\mat_mul/mult_37_G2/A1[5] ), .out(n3172) );
  inv U3878 ( .in(n3173), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[1].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[7] ) );
  inv U3879 ( .in(\mat_mul/mult_37_G2_G2_G1/A1[0] ), .out(n3174) );
  inv U3880 ( .in(n3175), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ) );
  inv U3881 ( .in(\mat_mul/mult_37_G2_G2_G1/A1[1] ), .out(n3176) );
  inv U3882 ( .in(n3177), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ) );
  inv U3883 ( .in(\mat_mul/mult_37_G2_G2_G1/A1[2] ), .out(n3178) );
  inv U3884 ( .in(n3179), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ) );
  inv U3885 ( .in(\mat_mul/mult_37_G2_G2_G1/A1[3] ), .out(n3180) );
  inv U3886 ( .in(n3181), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ) );
  inv U3887 ( .in(\mat_mul/mult_37_G2_G2_G1/A1[4] ), .out(n3182) );
  inv U3888 ( .in(n3183), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ) );
  inv U3889 ( .in(\mat_mul/mult_37_G2_G2_G1/A1[5] ), .out(n3184) );
  inv U3890 ( .in(n3185), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[7] ) );
  inv U3891 ( .in(\mat_mul/mult_37_G2_G1/A1[0] ), .out(n3186) );
  inv U3892 ( .in(n3187), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ) );
  inv U3893 ( .in(\mat_mul/mult_37_G2_G1/A1[1] ), .out(n3188) );
  inv U3894 ( .in(n3189), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[3] ) );
  inv U3895 ( .in(\mat_mul/mult_37_G2_G1/A1[2] ), .out(n3190) );
  inv U3896 ( .in(n3191), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ) );
  inv U3897 ( .in(\mat_mul/mult_37_G2_G1/A1[3] ), .out(n3192) );
  inv U3898 ( .in(n3193), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[5] ) );
  inv U3899 ( .in(\mat_mul/mult_37_G2_G1/A1[4] ), .out(n3194) );
  inv U3900 ( .in(n3195), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ) );
  inv U3901 ( .in(\mat_mul/mult_37_G2_G1/A1[5] ), .out(n3196) );
  inv U3902 ( .in(n3197), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[1].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[7] ) );
  inv U3903 ( .in(\mat_mul/mult_37_G2_G1_G1/A1[0] ), .out(n3198) );
  inv U3904 ( .in(n3199), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[2] ) );
  inv U3905 ( .in(\mat_mul/mult_37_G2_G1_G1/A1[1] ), .out(n3200) );
  inv U3906 ( .in(n3201), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[3] ) );
  inv U3907 ( .in(\mat_mul/mult_37_G2_G1_G1/A1[2] ), .out(n3202) );
  inv U3908 ( .in(n3203), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[4] ) );
  inv U3909 ( .in(\mat_mul/mult_37_G2_G1_G1/A1[3] ), .out(n3204) );
  inv U3910 ( .in(n3205), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[5] ) );
  inv U3911 ( .in(\mat_mul/mult_37_G2_G1_G1/A1[4] ), .out(n3206) );
  inv U3912 ( .in(n3207), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[6] ) );
  inv U3913 ( .in(\mat_mul/mult_37_G2_G1_G1/A1[5] ), .out(n3208) );
  inv U3914 ( .in(n3209), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[1].temp_res0_w[7] ) );
  inv U3915 ( .in(\mat_mul/mult_37/A1[0] ), .out(n3210) );
  inv U3916 ( .in(n3211), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[2] ) );
  inv U3917 ( .in(\mat_mul/mult_37/A1[1] ), .out(n3212) );
  inv U3918 ( .in(n3213), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[3] ) );
  inv U3919 ( .in(\mat_mul/mult_37/A1[2] ), .out(n3214) );
  inv U3920 ( .in(n3215), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[4] ) );
  inv U3921 ( .in(\mat_mul/mult_37/A1[3] ), .out(n3216) );
  inv U3922 ( .in(n3217), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[5] ) );
  inv U3923 ( .in(\mat_mul/mult_37/A1[4] ), .out(n3218) );
  inv U3924 ( .in(n3219), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[6] ) );
  inv U3925 ( .in(\mat_mul/mult_37/A1[5] ), .out(n3220) );
  inv U3926 ( .in(n3221), .out(
        \mat_mul/mul_mat_matrixproduct_wire_gen_block_1[0].mul_mat_matrixproduct_wire_gen_block_2[0].mul_mat_matrixproduct_wire_gen_block_3[0].temp_res0_w[7] ) );
  inv U3927 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/A1[0] ), .out(n3222) );
  inv U3928 ( .in(n3223), .out(m_kro[2]) );
  inv U3929 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/A1[1] ), .out(n3224) );
  inv U3930 ( .in(n3225), .out(m_kro[3]) );
  inv U3931 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/A1[2] ), .out(n3226) );
  inv U3932 ( .in(n3227), .out(m_kro[4]) );
  inv U3933 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/A1[3] ), .out(n3228) );
  inv U3934 ( .in(n3229), .out(m_kro[5]) );
  inv U3935 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/A1[4] ), .out(n3230) );
  inv U3936 ( .in(n3231), .out(m_kro[6]) );
  inv U3937 ( .in(\mat_kron/mult_40_G2_G2_G2_G2/A1[5] ), .out(n3232) );
  inv U3938 ( .in(n3233), .out(m_kro[7]) );
  inv U3939 ( .in(\mat_kron/mult_40_G2_G2_G2/A1[0] ), .out(n3234) );
  inv U3940 ( .in(n3235), .out(m_kro[10]) );
  inv U3941 ( .in(\mat_kron/mult_40_G2_G2_G2/A1[1] ), .out(n3236) );
  inv U3942 ( .in(n3237), .out(m_kro[11]) );
  inv U3943 ( .in(\mat_kron/mult_40_G2_G2_G2/A1[2] ), .out(n3238) );
  inv U3944 ( .in(n3239), .out(m_kro[12]) );
  inv U3945 ( .in(\mat_kron/mult_40_G2_G2_G2/A1[3] ), .out(n3240) );
  inv U3946 ( .in(n3241), .out(m_kro[13]) );
  inv U3947 ( .in(\mat_kron/mult_40_G2_G2_G2/A1[4] ), .out(n3242) );
  inv U3948 ( .in(n3243), .out(m_kro[14]) );
  inv U3949 ( .in(\mat_kron/mult_40_G2_G2_G2/A1[5] ), .out(n3244) );
  inv U3950 ( .in(n3245), .out(m_kro[15]) );
  inv U3951 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/A1[0] ), .out(n3246) );
  inv U3952 ( .in(n3247), .out(m_kro[34]) );
  inv U3953 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/A1[1] ), .out(n3248) );
  inv U3954 ( .in(n3249), .out(m_kro[35]) );
  inv U3955 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/A1[2] ), .out(n3250) );
  inv U3956 ( .in(n3251), .out(m_kro[36]) );
  inv U3957 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/A1[3] ), .out(n3252) );
  inv U3958 ( .in(n3253), .out(m_kro[37]) );
  inv U3959 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/A1[4] ), .out(n3254) );
  inv U3960 ( .in(n3255), .out(m_kro[38]) );
  inv U3961 ( .in(\mat_kron/mult_40_G2_G1_G2_G2/A1[5] ), .out(n3256) );
  inv U3962 ( .in(n3257), .out(m_kro[39]) );
  inv U3963 ( .in(\mat_kron/mult_40_G2_G2/A1[0] ), .out(n3258) );
  inv U3964 ( .in(n3259), .out(m_kro[42]) );
  inv U3965 ( .in(\mat_kron/mult_40_G2_G2/A1[1] ), .out(n3260) );
  inv U3966 ( .in(n3261), .out(m_kro[43]) );
  inv U3967 ( .in(\mat_kron/mult_40_G2_G2/A1[2] ), .out(n3262) );
  inv U3968 ( .in(n3263), .out(m_kro[44]) );
  inv U3969 ( .in(\mat_kron/mult_40_G2_G2/A1[3] ), .out(n3264) );
  inv U3970 ( .in(n3265), .out(m_kro[45]) );
  inv U3971 ( .in(\mat_kron/mult_40_G2_G2/A1[4] ), .out(n3266) );
  inv U3972 ( .in(n3267), .out(m_kro[46]) );
  inv U3973 ( .in(\mat_kron/mult_40_G2_G2/A1[5] ), .out(n3268) );
  inv U3974 ( .in(n3269), .out(m_kro[47]) );
  inv U3975 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/A1[0] ), .out(n3270) );
  inv U3976 ( .in(n3271), .out(m_kro[18]) );
  inv U3977 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/A1[1] ), .out(n3272) );
  inv U3978 ( .in(n3273), .out(m_kro[19]) );
  inv U3979 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/A1[2] ), .out(n3274) );
  inv U3980 ( .in(n3275), .out(m_kro[20]) );
  inv U3981 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/A1[3] ), .out(n3276) );
  inv U3982 ( .in(n3277), .out(m_kro[21]) );
  inv U3983 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/A1[4] ), .out(n3278) );
  inv U3984 ( .in(n3279), .out(m_kro[22]) );
  inv U3985 ( .in(\mat_kron/mult_40_G2_G2_G1_G2/A1[5] ), .out(n3280) );
  inv U3986 ( .in(n3281), .out(m_kro[23]) );
  inv U3987 ( .in(\mat_kron/mult_40_G2_G1_G2/A1[0] ), .out(n3282) );
  inv U3988 ( .in(n3283), .out(m_kro[26]) );
  inv U3989 ( .in(\mat_kron/mult_40_G2_G1_G2/A1[1] ), .out(n3284) );
  inv U3990 ( .in(n3285), .out(m_kro[27]) );
  inv U3991 ( .in(\mat_kron/mult_40_G2_G1_G2/A1[2] ), .out(n3286) );
  inv U3992 ( .in(n3287), .out(m_kro[28]) );
  inv U3993 ( .in(\mat_kron/mult_40_G2_G1_G2/A1[3] ), .out(n3288) );
  inv U3994 ( .in(n3289), .out(m_kro[29]) );
  inv U3995 ( .in(\mat_kron/mult_40_G2_G1_G2/A1[4] ), .out(n3290) );
  inv U3996 ( .in(n3291), .out(m_kro[30]) );
  inv U3997 ( .in(\mat_kron/mult_40_G2_G1_G2/A1[5] ), .out(n3292) );
  inv U3998 ( .in(n3293), .out(m_kro[31]) );
  inv U3999 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/A1[0] ), .out(n3294) );
  inv U4000 ( .in(n3295), .out(m_kro[50]) );
  inv U4001 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/A1[1] ), .out(n3296) );
  inv U4002 ( .in(n3297), .out(m_kro[51]) );
  inv U4003 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/A1[2] ), .out(n3298) );
  inv U4004 ( .in(n3299), .out(m_kro[52]) );
  inv U4005 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/A1[3] ), .out(n3300) );
  inv U4006 ( .in(n3301), .out(m_kro[53]) );
  inv U4007 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/A1[4] ), .out(n3302) );
  inv U4008 ( .in(n3303), .out(m_kro[54]) );
  inv U4009 ( .in(\mat_kron/mult_40_G2_G1_G1_G2/A1[5] ), .out(n3304) );
  inv U4010 ( .in(n3305), .out(m_kro[55]) );
  inv U4011 ( .in(\mat_kron/mult_40_G2/A1[0] ), .out(n3306) );
  inv U4012 ( .in(n3307), .out(m_kro[58]) );
  inv U4013 ( .in(\mat_kron/mult_40_G2/A1[1] ), .out(n3308) );
  inv U4014 ( .in(n3309), .out(m_kro[59]) );
  inv U4015 ( .in(\mat_kron/mult_40_G2/A1[2] ), .out(n3310) );
  inv U4016 ( .in(n3311), .out(m_kro[60]) );
  inv U4017 ( .in(\mat_kron/mult_40_G2/A1[3] ), .out(n3312) );
  inv U4018 ( .in(n3313), .out(m_kro[61]) );
  inv U4019 ( .in(\mat_kron/mult_40_G2/A1[4] ), .out(n3314) );
  inv U4020 ( .in(n3315), .out(m_kro[62]) );
  inv U4021 ( .in(\mat_kron/mult_40_G2/A1[5] ), .out(n3316) );
  inv U4022 ( .in(n3317), .out(m_kro[63]) );
  inv U4023 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/A1[0] ), .out(n3318) );
  inv U4024 ( .in(n3319), .out(m_kro[66]) );
  inv U4025 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/A1[1] ), .out(n3320) );
  inv U4026 ( .in(n3321), .out(m_kro[67]) );
  inv U4027 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/A1[2] ), .out(n3322) );
  inv U4028 ( .in(n3323), .out(m_kro[68]) );
  inv U4029 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/A1[3] ), .out(n3324) );
  inv U4030 ( .in(n3325), .out(m_kro[69]) );
  inv U4031 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/A1[4] ), .out(n3326) );
  inv U4032 ( .in(n3327), .out(m_kro[70]) );
  inv U4033 ( .in(\mat_kron/mult_40_G2_G2_G2_G1/A1[5] ), .out(n3328) );
  inv U4034 ( .in(n3329), .out(m_kro[71]) );
  inv U4035 ( .in(\mat_kron/mult_40_G2_G2_G1/A1[0] ), .out(n3330) );
  inv U4036 ( .in(n3331), .out(m_kro[74]) );
  inv U4037 ( .in(\mat_kron/mult_40_G2_G2_G1/A1[1] ), .out(n3332) );
  inv U4038 ( .in(n3333), .out(m_kro[75]) );
  inv U4039 ( .in(\mat_kron/mult_40_G2_G2_G1/A1[2] ), .out(n3334) );
  inv U4040 ( .in(n3335), .out(m_kro[76]) );
  inv U4041 ( .in(\mat_kron/mult_40_G2_G2_G1/A1[3] ), .out(n3336) );
  inv U4042 ( .in(n3337), .out(m_kro[77]) );
  inv U4043 ( .in(\mat_kron/mult_40_G2_G2_G1/A1[4] ), .out(n3338) );
  inv U4044 ( .in(n3339), .out(m_kro[78]) );
  inv U4045 ( .in(\mat_kron/mult_40_G2_G2_G1/A1[5] ), .out(n3340) );
  inv U4046 ( .in(n3341), .out(m_kro[79]) );
  inv U4047 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/A1[0] ), .out(n3342) );
  inv U4048 ( .in(n3343), .out(m_kro[98]) );
  inv U4049 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/A1[1] ), .out(n3344) );
  inv U4050 ( .in(n3345), .out(m_kro[99]) );
  inv U4051 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/A1[2] ), .out(n3346) );
  inv U4052 ( .in(n3347), .out(m_kro[100]) );
  inv U4053 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/A1[3] ), .out(n3348) );
  inv U4054 ( .in(n3349), .out(m_kro[101]) );
  inv U4055 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/A1[4] ), .out(n3350) );
  inv U4056 ( .in(n3351), .out(m_kro[102]) );
  inv U4057 ( .in(\mat_kron/mult_40_G2_G1_G2_G1/A1[5] ), .out(n3352) );
  inv U4058 ( .in(n3353), .out(m_kro[103]) );
  inv U4059 ( .in(\mat_kron/mult_40_G2_G1/A1[0] ), .out(n3354) );
  inv U4060 ( .in(n3355), .out(m_kro[106]) );
  inv U4061 ( .in(\mat_kron/mult_40_G2_G1/A1[1] ), .out(n3356) );
  inv U4062 ( .in(n3357), .out(m_kro[107]) );
  inv U4063 ( .in(\mat_kron/mult_40_G2_G1/A1[2] ), .out(n3358) );
  inv U4064 ( .in(n3359), .out(m_kro[108]) );
  inv U4065 ( .in(\mat_kron/mult_40_G2_G1/A1[3] ), .out(n3360) );
  inv U4066 ( .in(n3361), .out(m_kro[109]) );
  inv U4067 ( .in(\mat_kron/mult_40_G2_G1/A1[4] ), .out(n3362) );
  inv U4068 ( .in(n3363), .out(m_kro[110]) );
  inv U4069 ( .in(\mat_kron/mult_40_G2_G1/A1[5] ), .out(n3364) );
  inv U4070 ( .in(n3365), .out(m_kro[111]) );
  inv U4071 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/A1[0] ), .out(n3366) );
  inv U4072 ( .in(n3367), .out(m_kro[82]) );
  inv U4073 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/A1[1] ), .out(n3368) );
  inv U4074 ( .in(n3369), .out(m_kro[83]) );
  inv U4075 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/A1[2] ), .out(n3370) );
  inv U4076 ( .in(n3371), .out(m_kro[84]) );
  inv U4077 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/A1[3] ), .out(n3372) );
  inv U4078 ( .in(n3373), .out(m_kro[85]) );
  inv U4079 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/A1[4] ), .out(n3374) );
  inv U4080 ( .in(n3375), .out(m_kro[86]) );
  inv U4081 ( .in(\mat_kron/mult_40_G2_G2_G1_G1/A1[5] ), .out(n3376) );
  inv U4082 ( .in(n3377), .out(m_kro[87]) );
  inv U4083 ( .in(\mat_kron/mult_40_G2_G1_G1/A1[0] ), .out(n3378) );
  inv U4084 ( .in(n3379), .out(m_kro[90]) );
  inv U4085 ( .in(\mat_kron/mult_40_G2_G1_G1/A1[1] ), .out(n3380) );
  inv U4086 ( .in(n3381), .out(m_kro[91]) );
  inv U4087 ( .in(\mat_kron/mult_40_G2_G1_G1/A1[2] ), .out(n3382) );
  inv U4088 ( .in(n3383), .out(m_kro[92]) );
  inv U4089 ( .in(\mat_kron/mult_40_G2_G1_G1/A1[3] ), .out(n3384) );
  inv U4090 ( .in(n3385), .out(m_kro[93]) );
  inv U4091 ( .in(\mat_kron/mult_40_G2_G1_G1/A1[4] ), .out(n3386) );
  inv U4092 ( .in(n3387), .out(m_kro[94]) );
  inv U4093 ( .in(\mat_kron/mult_40_G2_G1_G1/A1[5] ), .out(n3388) );
  inv U4094 ( .in(n3389), .out(m_kro[95]) );
  inv U4095 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/A1[0] ), .out(n3390) );
  inv U4096 ( .in(n3391), .out(m_kro[114]) );
  inv U4097 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/A1[1] ), .out(n3392) );
  inv U4098 ( .in(n3393), .out(m_kro[115]) );
  inv U4099 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/A1[2] ), .out(n3394) );
  inv U4100 ( .in(n3395), .out(m_kro[116]) );
  inv U4101 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/A1[3] ), .out(n3396) );
  inv U4102 ( .in(n3397), .out(m_kro[117]) );
  inv U4103 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/A1[4] ), .out(n3398) );
  inv U4104 ( .in(n3399), .out(m_kro[118]) );
  inv U4105 ( .in(\mat_kron/mult_40_G2_G1_G1_G1/A1[5] ), .out(n3400) );
  inv U4106 ( .in(n3401), .out(m_kro[119]) );
  inv U4107 ( .in(\mat_kron/mult_40/A1[0] ), .out(n3402) );
  inv U4108 ( .in(n3403), .out(m_kro[122]) );
  inv U4109 ( .in(\mat_kron/mult_40/A1[1] ), .out(n3404) );
  inv U4110 ( .in(n3405), .out(m_kro[123]) );
  inv U4111 ( .in(\mat_kron/mult_40/A1[2] ), .out(n3406) );
  inv U4112 ( .in(n3407), .out(m_kro[124]) );
  inv U4113 ( .in(\mat_kron/mult_40/A1[3] ), .out(n3408) );
  inv U4114 ( .in(n3409), .out(m_kro[125]) );
  inv U4115 ( .in(\mat_kron/mult_40/A1[4] ), .out(n3410) );
  inv U4116 ( .in(n3411), .out(m_kro[126]) );
  inv U4117 ( .in(\mat_kron/mult_40/A1[5] ), .out(n3412) );
  inv U4118 ( .in(n3413), .out(m_kro[127]) );
endmodule



